LIBRARY ieee;
USE ieee.STD_LOGIC_1164.ALL;

PACKAGE constants_pkg IS
    CONSTANT DATAWIDTH    : INTEGER := 13;
    CONSTANT ADDRWIDTH    : INTEGER := 12;
    CONSTANT SAMPLINGFREQ : INTEGER := 6249;
END PACKAGE;