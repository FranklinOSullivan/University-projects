LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY power_signal_rom IS
    PORT (
        clk : IN STD_LOGIC;
        address : IN INTEGER RANGE 0 TO 1599; -- 10 cycles * 16000 samples/s / 50 Hz
        data_out : OUT unsigned(15 DOWNTO 0) -- 8-bit output
    );
END power_signal_rom;

ARCHITECTURE Behavioral OF power_signal_rom IS
    TYPE rom_type IS ARRAY (0 TO 1599) OF unsigned(15 DOWNTO 0);
    ---FAT array with 1600 samples of the power signal
    SIGNAL rom : rom_type := (
        0 => "1110110111010000",
        1 => "1111001110010000",
        2 => "1111011110100000",
        3 => "1111101101000000",
        4 => "1110100111000000",
        5 => "1111010011000000",
        6 => "1111010000000000",
        7 => "1111000101110000",
        8 => "1110011010000000",
        9 => "1110101100010000",
        10 => "1101111000100000",
        11 => "1101110110110000",
        12 => "1101011111110000",
        13 => "1101011001000000",
        14 => "1100111101110000",
        15 => "1101000011100000",
        16 => "1100000101010000",
        17 => "1011010010010000",
        18 => "1100000011000000",
        19 => "1011100001110000",
        20 => "1001110000110000",
        21 => "1010111100100000",
        22 => "1001110010000000",
        23 => "1001111000110000",
        24 => "1001010011010000",
        25 => "1000101110010000",
        26 => "1000011010110000",
        27 => "0111110011010000",
        28 => "0111000101010000",
        29 => "0111010100010000",
        30 => "0111001000010000",
        31 => "0110100110010000",
        32 => "0111001100110000",
        33 => "0101110011100000",
        34 => "0110000000010000",
        35 => "0110010011000000",
        36 => "0101101100000000",
        37 => "0101001010000000",
        38 => "0101110111000000",
        39 => "0101110101100000",
        40 => "0100010110000000",
        41 => "0100000111110000",
        42 => "0101000100100000",
        43 => "0100111110110000",
        44 => "0101100111000000",
        45 => "0100011110010000",
        46 => "0100101001100000",
        47 => "0100011100010000",
        48 => "0100001001010000",
        49 => "0100110000010000",
        50 => "0011111111010000",
        51 => "0100101111110000",
        52 => "0100000010110000",
        53 => "0011110000100000",
        54 => "0011011011010000",
        55 => "0011101011110000",
        56 => "0011101111100000",
        57 => "0100000100100000",
        58 => "0010010001010000",
        59 => "0011010010000000",
        60 => "0011100000110000",
        61 => "0010101010010000",
        62 => "0010001010110000",
        63 => "0010001111000000",
        64 => "0011100111010000",
        65 => "0010011011100000",
        66 => "0011001100010000",
        67 => "0010010011010000",
        68 => "0010111110110000",
        69 => "0010111000110000",
        70 => "0010101011110000",
        71 => "0011000001010000",
        72 => "0011011001000000",
        73 => "0010000000010000",
        74 => "0010101101010000",
        75 => "0010011100000000",
        76 => "0010100100000000",
        77 => "0001111111000000",
        78 => "0001111000000000",
        79 => "0010101101110000",
        80 => "0001110101110000",
        81 => "0010011011000000",
        82 => "0010011000000000",
        83 => "0001111111010000",
        84 => "0010100101110000",
        85 => "0001101110100000",
        86 => "0010011111100000",
        87 => "0010101110110000",
        88 => "0010010110010000",
        89 => "0010001001110000",
        90 => "0010001010110000",
        91 => "0001100111100000",
        92 => "0010100000010000",
        93 => "0001111000000000",
        94 => "0010110110000000",
        95 => "0010001111100000",
        96 => "0010001100010000",
        97 => "0010101101010000",
        98 => "0010111001010000",
        99 => "0010000010000000",
        100 => "0010101100100000",
        101 => "0010011011000000",
        102 => "0010101000100000",
        103 => "0010001010100000",
        104 => "0010100011110000",
        105 => "0010110000000000",
        106 => "0011100111100000",
        107 => "0010011000000000",
        108 => "0010101101110000",
        109 => "0011000111000000",
        110 => "0010110010010000",
        111 => "0011100010110000",
        112 => "0011011111000000",
        113 => "0011000010110000",
        114 => "0011011110010000",
        115 => "0011110000100000",
        116 => "0011000011110000",
        117 => "0010101010000000",
        118 => "0010110000100000",
        119 => "0010110110000000",
        120 => "0010101000010000",
        121 => "0010111010000000",
        122 => "0010110010010000",
        123 => "0011011011110000",
        124 => "0011110100010000",
        125 => "0011100010010000",
        126 => "0011101001110000",
        127 => "0010111101110000",
        128 => "0010111010000000",
        129 => "0010110000000000",
        130 => "0010100110110000",
        131 => "0011100101110000",
        132 => "0100001000100000",
        133 => "0011001000110000",
        134 => "0011111010010000",
        135 => "0010101111000000",
        136 => "0011110111010000",
        137 => "0100001110010000",
        138 => "0011010000000000",
        139 => "0011100101100000",
        140 => "0010110010000000",
        141 => "0011000101000000",
        142 => "0011101111110000",
        143 => "0011011110100000",
        144 => "0011101100110000",
        145 => "0010111110110000",
        146 => "0011001001100000",
        147 => "0011000110110000",
        148 => "0010001100100000",
        149 => "0010110011110000",
        150 => "0011000101110000",
        151 => "0010010100100000",
        152 => "0010000010110000",
        153 => "0001100000100000",
        154 => "0001110010000000",
        155 => "0001110011110000",
        156 => "0001000101110000",
        157 => "0010011000110000",
        158 => "0001011010100000",
        159 => "0001110011100000",
        160 => "0001000101000000",
        161 => "0001010001010000",
        162 => "0000110010100000",
        163 => "0001011000110000",
        164 => "0000101001110000",
        165 => "0001001111100000",
        166 => "0000001011000000",
        167 => "0000110100100000",
        168 => "0001000010010000",
        169 => "0001110100010000",
        170 => "0010010001110000",
        171 => "0001100010000000",
        172 => "0001101100100000",
        173 => "0010010001010000",
        174 => "0010101010110000",
        175 => "0010110100110000",
        176 => "0011001010010000",
        177 => "0100001011000000",
        178 => "0100010000010000",
        179 => "0100100111010000",
        180 => "0100010110100000",
        181 => "0101100000100000",
        182 => "0101010111110000",
        183 => "0101110100110000",
        184 => "0110110001100000",
        185 => "0111011001000000",
        186 => "0111011000010000",
        187 => "0111110101100000",
        188 => "0111111000000000",
        189 => "1000110100000000",
        190 => "1000100011110000",
        191 => "1000100011010000",
        192 => "1000001011000000",
        193 => "1001101001000000",
        194 => "1001110100110000",
        195 => "1001101100100000",
        196 => "1001011011000000",
        197 => "1010111110100000",
        198 => "1010101101000000",
        199 => "1010011100000000",
        200 => "1011011010110000",
        201 => "1010000111100000",
        202 => "1011000010000000",
        203 => "1011110111110000",
        204 => "1011010101000000",
        205 => "1010111100010000",
        206 => "1011001010110000",
        207 => "1011001010000000",
        208 => "1011001100100000",
        209 => "1011101010110000",
        210 => "1011001111000000",
        211 => "1011101011000000",
        212 => "1100000111110000",
        213 => "1100000100110000",
        214 => "1011010000110000",
        215 => "1100100000100000",
        216 => "1011111111010000",
        217 => "1100011111110000",
        218 => "1100101000110000",
        219 => "1101001011010000",
        220 => "1100110001100000",
        221 => "1011111000010000",
        222 => "1100000100000000",
        223 => "1101110000110000",
        224 => "1101000100000000",
        225 => "1100111101100000",
        226 => "1101000000100000",
        227 => "1101001101000000",
        228 => "1101000010100000",
        229 => "1100110100100000",
        230 => "1100111001110000",
        231 => "1101010000010000",
        232 => "1100110110110000",
        233 => "1101101010000000",
        234 => "1101011011000000",
        235 => "1100111011110000",
        236 => "1100110001010000",
        237 => "1100101000010000",
        238 => "1101010110100000",
        239 => "1101100000000000",
        240 => "1101010100110000",
        241 => "1110000110110000",
        242 => "1101001010000000",
        243 => "1100111011100000",
        244 => "1101111011100000",
        245 => "1101011001010000",
        246 => "1100110111010000",
        247 => "1100100100110000",
        248 => "1101111011000000",
        249 => "1101110110010000",
        250 => "1101111010100000",
        251 => "1101011101000000",
        252 => "1101010100110000",
        253 => "1101111101000000",
        254 => "1101110110100000",
        255 => "1101101011010000",
        256 => "1101101001010000",
        257 => "1101100100010000",
        258 => "1101011101000000",
        259 => "1101011111110000",
        260 => "1110011111000000",
        261 => "1101011111010000",
        262 => "1110000011010000",
        263 => "1101110111010000",
        264 => "1101110011000000",
        265 => "1101110011010000",
        266 => "1101011110110000",
        267 => "1110001110010000",
        268 => "1100110000110000",
        269 => "1100001001000000",
        270 => "1101010000110000",
        271 => "1100010100110000",
        272 => "1100111100010000",
        273 => "1101001110110000",
        274 => "1101100011110000",
        275 => "1100100001000000",
        276 => "1101010010100000",
        277 => "1101000001010000",
        278 => "1100100100100000",
        279 => "1101010011110000",
        280 => "1100100110100000",
        281 => "1101001111000000",
        282 => "1100100001000000",
        283 => "1100110000100000",
        284 => "1100111110110000",
        285 => "1101100111010000",
        286 => "1101010001000000",
        287 => "1100101101010000",
        288 => "1101001110010000",
        289 => "1100100110100000",
        290 => "1101010101100000",
        291 => "1100100001000000",
        292 => "1011110010010000",
        293 => "1100000011100000",
        294 => "1100000010100000",
        295 => "1100001001110000",
        296 => "1101010011010000",
        297 => "1101001001000000",
        298 => "1101000110000000",
        299 => "1100100111000000",
        300 => "1101000110110000",
        301 => "1101010000010000",
        302 => "1100010001010000",
        303 => "1100001010010000",
        304 => "1011111000100000",
        305 => "1100000101100000",
        306 => "1101100101100000",
        307 => "1100101000000000",
        308 => "1100101101110000",
        309 => "1101011011010000",
        310 => "1100100010110000",
        311 => "1100110110110000",
        312 => "1100110111110000",
        313 => "1110011101010000",
        314 => "1101110010100000",
        315 => "1110011101000000",
        316 => "1110101001110000",
        317 => "1110011110100000",
        318 => "1110110001100000",
        319 => "1110100011100000",
        320 => "1111101111000000",
        321 => "1110111010010000",
        322 => "1110010010110000",
        323 => "1111110011110000",
        324 => "1110100101010000",
        325 => "1110001100010000",
        326 => "1110100100000000",
        327 => "1111000000100000",
        328 => "1110011110010000",
        329 => "1110001011010000",
        330 => "1110010000100000",
        331 => "1110100101000000",
        332 => "1101110111100000",
        333 => "1101100110010000",
        334 => "1101001001100000",
        335 => "1101000000100000",
        336 => "1100011011010000",
        337 => "1011001011000000",
        338 => "1100100111000000",
        339 => "1011111000100000",
        340 => "1010100110110000",
        341 => "1001010100000000",
        342 => "1001111010110000",
        343 => "1001001110110000",
        344 => "1000101111110000",
        345 => "0111111001000000",
        346 => "0111011111010000",
        347 => "0111100010100000",
        348 => "0111101100000000",
        349 => "0111110000100000",
        350 => "0110111100110000",
        351 => "0110111101010000",
        352 => "0110100101100000",
        353 => "0110110100110000",
        354 => "0101111111010000",
        355 => "0101110011110000",
        356 => "0101100010000000",
        357 => "0101000010100000",
        358 => "0101100010010000",
        359 => "0100100000110000",
        360 => "0101101100000000",
        361 => "0101010011000000",
        362 => "0101001101100000",
        363 => "0100100010010000",
        364 => "0100110001110000",
        365 => "0101000010110000",
        366 => "0100010011100000",
        367 => "0011111100000000",
        368 => "0100111011110000",
        369 => "0011101100010000",
        370 => "0100100010110000",
        371 => "0100000101000000",
        372 => "0100010111110000",
        373 => "0011110110110000",
        374 => "0100001000000000",
        375 => "0011010001010000",
        376 => "0011010000000000",
        377 => "0011011101000000",
        378 => "0010101011000000",
        379 => "0011110001110000",
        380 => "0011011010000000",
        381 => "0010101110000000",
        382 => "0011001000110000",
        383 => "0010010000000000",
        384 => "0010011001010000",
        385 => "0010111111100000",
        386 => "0011000000100000",
        387 => "0010101111000000",
        388 => "0010100111000000",
        389 => "0010010001000000",
        390 => "0011001000000000",
        391 => "0010101011010000",
        392 => "0010001000010000",
        393 => "0010111011100000",
        394 => "0010100011000000",
        395 => "0011100100010000",
        396 => "0011011000010000",
        397 => "0010001111100000",
        398 => "0011010101100000",
        399 => "0010100011110000",
        400 => "0001110010110000",
        401 => "0001110001010000",
        402 => "0010001101100000",
        403 => "0010010000100000",
        404 => "0010110000100000",
        405 => "0011011110100000",
        406 => "0010100011000000",
        407 => "0010011101000000",
        408 => "0010001011000000",
        409 => "0010010100110000",
        410 => "0010111011010000",
        411 => "0011001101010000",
        412 => "0010000010110000",
        413 => "0010100001000000",
        414 => "0010000100000000",
        415 => "0010100100010000",
        416 => "0010011101100000",
        417 => "0010110000110000",
        418 => "0010100101110000",
        419 => "0010000101110000",
        420 => "0010100001110000",
        421 => "0010010111110000",
        422 => "0011010000000000",
        423 => "0010110001110000",
        424 => "0010000000000000",
        425 => "0011001010100000",
        426 => "0011010101010000",
        427 => "0011001011110000",
        428 => "0010011011100000",
        429 => "0010100001110000",
        430 => "0010000111000000",
        431 => "0010001011000000",
        432 => "0010100110010000",
        433 => "0011000101100000",
        434 => "0010011111100000",
        435 => "0011111010100000",
        436 => "0011010011010000",
        437 => "0011000101010000",
        438 => "0010101100110000",
        439 => "0011110110110000",
        440 => "0010110011010000",
        441 => "0011010011100000",
        442 => "0010111000110000",
        443 => "0010101010110000",
        444 => "0010001101110000",
        445 => "0011001100000000",
        446 => "0011111010100000",
        447 => "0010010010110000",
        448 => "0010110110010000",
        449 => "0010011011010000",
        450 => "0011110110010000",
        451 => "0011100010000000",
        452 => "0010011010110000",
        453 => "0010100111010000",
        454 => "0010111111110000",
        455 => "0011010110110000",
        456 => "0010011111110000",
        457 => "0010110000110000",
        458 => "0010110000110000",
        459 => "0010101100000000",
        460 => "0011111101000000",
        461 => "0011001011010000",
        462 => "0011110010010000",
        463 => "0010111110000000",
        464 => "0010111101110000",
        465 => "0010111011010000",
        466 => "0011011011000000",
        467 => "0010101100100000",
        468 => "0001111111000000",
        469 => "0010000101000000",
        470 => "0001111101000000",
        471 => "0010011110010000",
        472 => "0010010010000000",
        473 => "0010000101000000",
        474 => "0001001111000000",
        475 => "0010000010110000",
        476 => "0001010010010000",
        477 => "0001000010000000",
        478 => "0001110101100000",
        479 => "0000011111110000",
        480 => "0000001001110000",
        481 => "0000001011100000",
        482 => "0001010010110000",
        483 => "0000100001100000",
        484 => "0000011101000000",
        485 => "0000110100000000",
        486 => "0001000010010000",
        487 => "0000100001000000",
        488 => "0000111110000000",
        489 => "0001000001010000",
        490 => "0001111101000000",
        491 => "0010100011000000",
        492 => "0001011100010000",
        493 => "0010001110100000",
        494 => "0001111101100000",
        495 => "0011001100010000",
        496 => "0010110110100000",
        497 => "0100010111010000",
        498 => "0011111010110000",
        499 => "0100001110000000",
        500 => "0101101011100000",
        501 => "0101101000000000",
        502 => "0110000110000000",
        503 => "0110101101010000",
        504 => "0111011110110000",
        505 => "0111010110110000",
        506 => "1000001111000000",
        507 => "0111011100100000",
        508 => "1000110010100000",
        509 => "1000000011100000",
        510 => "1001110101110000",
        511 => "1001010110100000",
        512 => "1001110011000000",
        513 => "1001100001100000",
        514 => "1010010010000000",
        515 => "1001011111110000",
        516 => "1010010110100000",
        517 => "1001101101000000",
        518 => "1010001101110000",
        519 => "1010010111000000",
        520 => "1010010000010000",
        521 => "1010100010110000",
        522 => "1010100101000000",
        523 => "1010100101010000",
        524 => "1010101101110000",
        525 => "1011000100000000",
        526 => "1011011010110000",
        527 => "1011001011100000",
        528 => "1011010100010000",
        529 => "1011010011100000",
        530 => "1011011100100000",
        531 => "1011111100000000",
        532 => "1011100101100000",
        533 => "1011111111000000",
        534 => "1100000101000000",
        535 => "1011110110010000",
        536 => "1011101101100000",
        537 => "1011101000110000",
        538 => "1100011110000000",
        539 => "1100100110100000",
        540 => "1100001010110000",
        541 => "1100101010000000",
        542 => "1101000011110000",
        543 => "1101010100100000",
        544 => "1100011110010000",
        545 => "1101000100100000",
        546 => "1100110000110000",
        547 => "1101000101100000",
        548 => "1101110000100000",
        549 => "1101100011110000",
        550 => "1100100110010000",
        551 => "1101001011010000",
        552 => "1101101000110000",
        553 => "1100110011000000",
        554 => "1101110111100000",
        555 => "1101010100110000",
        556 => "1101011111000000",
        557 => "1101101011010000",
        558 => "1101101110000000",
        559 => "1101011100100000",
        560 => "1101100000100000",
        561 => "1101110110100000",
        562 => "1101000110010000",
        563 => "1110000100100000",
        564 => "1101010011110000",
        565 => "1101001001110000",
        566 => "1101011110010000",
        567 => "1100110101100000",
        568 => "1101011010010000",
        569 => "1101110000010000",
        570 => "1101011100010000",
        571 => "1110001000000000",
        572 => "1101010001110000",
        573 => "1101001001010000",
        574 => "1101100110100000",
        575 => "1110000000110000",
        576 => "1101100111010000",
        577 => "1101111101010000",
        578 => "1101000110000000",
        579 => "1100111011100000",
        580 => "1101100101110000",
        581 => "1100100000100000",
        582 => "1101011111000000",
        583 => "1100110100010000",
        584 => "1100111100100000",
        585 => "1101001100110000",
        586 => "1101011110000000",
        587 => "1101010000010000",
        588 => "1100111000100000",
        589 => "1101011001010000",
        590 => "1101101000100000",
        591 => "1100011110110000",
        592 => "1100101100100000",
        593 => "1100111110010000",
        594 => "1100111101110000",
        595 => "1100110010010000",
        596 => "1101001010110000",
        597 => "1101000001100000",
        598 => "1100101101010000",
        599 => "1100111000000000",
        600 => "1100100000100000",
        601 => "1100011110000000",
        602 => "1100111101010000",
        603 => "1101110100110000",
        604 => "1101101100100000",
        605 => "1100110110010000",
        606 => "1100111100000000",
        607 => "1100001010010000",
        608 => "1101000111110000",
        609 => "1100100101100000",
        610 => "1101010101110000",
        611 => "1100001101110000",
        612 => "1101000011100000",
        613 => "1100110101000000",
        614 => "1100111100000000",
        615 => "1100000010000000",
        616 => "1011111011100000",
        617 => "1101001010010000",
        618 => "1011110111010000",
        619 => "1101010111110000",
        620 => "1100010000000000",
        621 => "1100010110010000",
        622 => "1101010111000000",
        623 => "1101000010100000",
        624 => "1101010100110000",
        625 => "1100110011100000",
        626 => "1100110110000000",
        627 => "1100101110010000",
        628 => "1101110101100000",
        629 => "1101000001000000",
        630 => "1100110111110000",
        631 => "1101110111110000",
        632 => "1100100100100000",
        633 => "1101110101000000",
        634 => "1110000001010000",
        635 => "1110011000010000",
        636 => "1110101010110000",
        637 => "1110101011010000",
        638 => "1110100101100000",
        639 => "1110100111000000",
        640 => "1111110100100000",
        641 => "1111001010110000",
        642 => "1101111100000000",
        643 => "1101111111100000",
        644 => "1111001101010000",
        645 => "1110101100010000",
        646 => "1110110000100000",
        647 => "1111001001000000",
        648 => "1110100110000000",
        649 => "1101111100000000",
        650 => "1101101111000000",
        651 => "1110010010000000",
        652 => "1101011010110000",
        653 => "1100111011010000",
        654 => "1011111001100000",
        655 => "1100111111000000",
        656 => "1100001011000000",
        657 => "1100000010000000",
        658 => "1010000110010000",
        659 => "1011000011010000",
        660 => "1010101110000000",
        661 => "1001101100110000",
        662 => "1010010101010000",
        663 => "1000101101010000",
        664 => "1001111010010000",
        665 => "1000100101000000",
        666 => "0111100110000000",
        667 => "1000100010110000",
        668 => "0111001000100000",
        669 => "0111010010000000",
        670 => "0111011000010000",
        671 => "0110111101110000",
        672 => "0110010011000000",
        673 => "0111001010100000",
        674 => "0110011100000000",
        675 => "0101000011100000",
        676 => "0101010001100000",
        677 => "0100110101110000",
        678 => "0101110111100000",
        679 => "0100110011000000",
        680 => "0100101000110000",
        681 => "0100111101100000",
        682 => "0101001111000000",
        683 => "0101010101000000",
        684 => "0011110100100000",
        685 => "0100101101000000",
        686 => "0100100011010000",
        687 => "0100011010110000",
        688 => "0011111110000000",
        689 => "0011111011110000",
        690 => "0011101101100000",
        691 => "0100011100100000",
        692 => "0011110100110000",
        693 => "0011011001000000",
        694 => "0011101001100000",
        695 => "0011111111100000",
        696 => "0011010100110000",
        697 => "0011100011000000",
        698 => "0010110011100000",
        699 => "0011110100000000",
        700 => "0011100110000000",
        701 => "0011100011100000",
        702 => "0011000010000000",
        703 => "0011010000010000",
        704 => "0011100100000000",
        705 => "0001110111010000",
        706 => "0011010110000000",
        707 => "0010110111100000",
        708 => "0011001111000000",
        709 => "0010101111010000",
        710 => "0010101100000000",
        711 => "0010111001100000",
        712 => "0010110011110000",
        713 => "0010100001110000",
        714 => "0010001000000000",
        715 => "0010000000100000",
        716 => "0011000000100000",
        717 => "0010111000110000",
        718 => "0011001010100000",
        719 => "0010001000110000",
        720 => "0010111110110000",
        721 => "0010101100010000",
        722 => "0010101100110000",
        723 => "0010010001010000",
        724 => "0010010011110000",
        725 => "0010100111100000",
        726 => "0011001000110000",
        727 => "0010001100010000",
        728 => "0010010101110000",
        729 => "0001110101110000",
        730 => "0010000110110000",
        731 => "0001111100100000",
        732 => "0010001010100000",
        733 => "0010010111100000",
        734 => "0001111101000000",
        735 => "0010011110000000",
        736 => "0010001111100000",
        737 => "0010110110110000",
        738 => "0010000010110000",
        739 => "0010100100100000",
        740 => "0001100111010000",
        741 => "0001010111110000",
        742 => "0010101110110000",
        743 => "0011001001110000",
        744 => "0010001010110000",
        745 => "0010101101100000",
        746 => "0100011111010000",
        747 => "0010100100100000",
        748 => "0010111001000000",
        749 => "0010111010100000",
        750 => "0010100111000000",
        751 => "0010101011000000",
        752 => "0011011001110000",
        753 => "0011100011010000",
        754 => "0010011100110000",
        755 => "0010110010000000",
        756 => "0011010010010000",
        757 => "0010111111000000",
        758 => "0010011100110000",
        759 => "0011010001110000",
        760 => "0010111010110000",
        761 => "0010001011110000",
        762 => "0010111000000000",
        763 => "0010110000010000",
        764 => "0010101100100000",
        765 => "0010111011010000",
        766 => "0010100010010000",
        767 => "0011001110100000",
        768 => "0011100100100000",
        769 => "0011111100000000",
        770 => "0010110000010000",
        771 => "0011100111100000",
        772 => "0100011010000000",
        773 => "0011100101000000",
        774 => "0011011110000000",
        775 => "0010110011010000",
        776 => "0010111100010000",
        777 => "0011001000110000",
        778 => "0011001011000000",
        779 => "0011001011000000",
        780 => "0010101001100000",
        781 => "0010011100110000",
        782 => "0010100001110000",
        783 => "0011000010000000",
        784 => "0011011101010000",
        785 => "0011000001110000",
        786 => "0011100101010000",
        787 => "0010001101100000",
        788 => "0010001110000000",
        789 => "0010110010110000",
        790 => "0010101100110000",
        791 => "0010010110100000",
        792 => "0001101010110000",
        793 => "0001001110100000",
        794 => "0001101100100000",
        795 => "0001000000110000",
        796 => "0001101011110000",
        797 => "0001110110110000",
        798 => "0000001001110000",
        799 => "0001001011100000",
        800 => "0000110101110000",
        801 => "0000100111010000",
        802 => "0000101011000000",
        803 => "0001010000100000",
        804 => "0000110100100000",
        805 => "0000111011000000",
        806 => "0001000011110000",
        807 => "0000110100000000",
        808 => "0001000110010000",
        809 => "0001110110000000",
        810 => "0010000101100000",
        811 => "0010000111010000",
        812 => "0010010000110000",
        813 => "0010110100110000",
        814 => "0011001110110000",
        815 => "0011101100000000",
        816 => "0011011011100000",
        817 => "0100100000000000",
        818 => "0101010100100000",
        819 => "0100000100010000",
        820 => "0110000100000000",
        821 => "0101001010010000",
        822 => "0110000111110000",
        823 => "0110110011100000",
        824 => "0111000110010000",
        825 => "0110110100000000",
        826 => "0110011000110000",
        827 => "0111110000010000",
        828 => "0111111010000000",
        829 => "1001001010010000",
        830 => "1000110010010000",
        831 => "1000110010110000",
        832 => "1001101001000000",
        833 => "1001011100110000",
        834 => "1001101100010000",
        835 => "1001001100110000",
        836 => "1010001001010000",
        837 => "1010010101100000",
        838 => "1010001001100000",
        839 => "1010100011100000",
        840 => "1011001010110000",
        841 => "1010101000000000",
        842 => "1010111111100000",
        843 => "1010110101110000",
        844 => "1010110001110000",
        845 => "1011000000100000",
        846 => "1011001001100000",
        847 => "1011000001110000",
        848 => "1011100110000000",
        849 => "1100000001000000",
        850 => "1100001011110000",
        851 => "1011111100010000",
        852 => "1011111011010000",
        853 => "1011101011110000",
        854 => "1100110100100000",
        855 => "1100101111000000",
        856 => "1100110011110000",
        857 => "1100100011000000",
        858 => "1100110010110000",
        859 => "1100101000100000",
        860 => "1100011011000000",
        861 => "1101001011000000",
        862 => "1100011001110000",
        863 => "1100110000010000",
        864 => "1101100000010000",
        865 => "1100101001110000",
        866 => "1101010011100000",
        867 => "1100010001010000",
        868 => "1101010001000000",
        869 => "1101101010000000",
        870 => "1101001001000000",
        871 => "1101001000010000",
        872 => "1100111110010000",
        873 => "1101100100110000",
        874 => "1101001011110000",
        875 => "1100111100100000",
        876 => "1101010001000000",
        877 => "1101001101100000",
        878 => "1101010100110000",
        879 => "1101100000000000",
        880 => "1101100010100000",
        881 => "1101010100010000",
        882 => "1110000001100000",
        883 => "1101110100010000",
        884 => "1101110101010000",
        885 => "1100111001110000",
        886 => "1101010010100000",
        887 => "1101011101100000",
        888 => "1101011110010000",
        889 => "1101100010110000",
        890 => "1101011100110000",
        891 => "1101101011010000",
        892 => "1101001011000000",
        893 => "1100101110000000",
        894 => "1101110101010000",
        895 => "1101101100010000",
        896 => "1110000011000000",
        897 => "1100110011100000",
        898 => "1101101001000000",
        899 => "1101010101000000",
        900 => "1101100010010000",
        901 => "1101011101100000",
        902 => "1101010101110000",
        903 => "1101101010000000",
        904 => "1100111111000000",
        905 => "1100111110000000",
        906 => "1101100000000000",
        907 => "1101000110100000",
        908 => "1100010111100000",
        909 => "1101000011000000",
        910 => "1100011100000000",
        911 => "1101001101010000",
        912 => "1100011000010000",
        913 => "1100111001000000",
        914 => "1100100101000000",
        915 => "1100101011110000",
        916 => "1101101000100000",
        917 => "1100100000000000",
        918 => "1100111001110000",
        919 => "1100110101010000",
        920 => "1100110010010000",
        921 => "1100111011010000",
        922 => "1100101000110000",
        923 => "1100001111110000",
        924 => "1100011110100000",
        925 => "1101101110010000",
        926 => "1100011110010000",
        927 => "1101101101100000",
        928 => "1100110100000000",
        929 => "1100111111100000",
        930 => "1100010100010000",
        931 => "1101000001110000",
        932 => "1101011101100000",
        933 => "1100101001010000",
        934 => "1011111010010000",
        935 => "1101011110100000",
        936 => "1101000100010000",
        937 => "1100101111110000",
        938 => "1100011111000000",
        939 => "1101010000000000",
        940 => "1100100110100000",
        941 => "1101001000110000",
        942 => "1100011011010000",
        943 => "1100010011100000",
        944 => "1101011111000000",
        945 => "1100101011000000",
        946 => "1100111000000000",
        947 => "1100010101000000",
        948 => "1101010110010000",
        949 => "1101011011110000",
        950 => "1101111111000000",
        951 => "1101001100110000",
        952 => "1110001111100000",
        953 => "1110000101100000",
        954 => "1110000111010000",
        955 => "1110011111110000",
        956 => "1110000100100000",
        957 => "1111011111010000",
        958 => "1110010111100000",
        959 => "1110101110100000",
        960 => "1111011100000000",
        961 => "1111011010110000",
        962 => "1110101110100000",
        963 => "1111111111110000",
        964 => "1110101001100000",
        965 => "1110110110000000",
        966 => "1110111010000000",
        967 => "1111011100110000",
        968 => "1110010000000000",
        969 => "1110000010000000",
        970 => "1101101111100000",
        971 => "1110011100110000",
        972 => "1101110001010000",
        973 => "1100101110000000",
        974 => "1101100000000000",
        975 => "1100001110010000",
        976 => "1100100010100000",
        977 => "1011111010110000",
        978 => "1011001101000000",
        979 => "1010111001110000",
        980 => "1010110111000000",
        981 => "1010010010100000",
        982 => "1001010000000000",
        983 => "1001011100010000",
        984 => "1000011010010000",
        985 => "1000011101010000",
        986 => "1000001010000000",
        987 => "0111100100100000",
        988 => "0111001011100000",
        989 => "0111001010000000",
        990 => "0111010111110000",
        991 => "0110100100100000",
        992 => "0110011101000000",
        993 => "0101110101100000",
        994 => "0110010000010000",
        995 => "0101100000010000",
        996 => "0101110111010000",
        997 => "0110000101010000",
        998 => "0100110110110000",
        999 => "0101101100000000",
        1000 => "0100110000110000",
        1001 => "0100011000110000",
        1002 => "0100010000000000",
        1003 => "0101011011010000",
        1004 => "0100100100110000",
        1005 => "0100010000110000",
        1006 => "0100110100000000",
        1007 => "0101000011110000",
        1008 => "0101000011110000",
        1009 => "0100001011000000",
        1010 => "0101010001100000",
        1011 => "0100001101000000",
        1012 => "0100101000100000",
        1013 => "0011100010100000",
        1014 => "0011101110000000",
        1015 => "0011101011100000",
        1016 => "0011001110110000",
        1017 => "0011010001000000",
        1018 => "0011001101110000",
        1019 => "0011100011110000",
        1020 => "0011100010110000",
        1021 => "0010110010100000",
        1022 => "0010101101000000",
        1023 => "0011001110010000",
        1024 => "0010011000110000",
        1025 => "0010110001110000",
        1026 => "0011100000010000",
        1027 => "0011000001010000",
        1028 => "0011011000010000",
        1029 => "0001110011000000",
        1030 => "0010001100100000",
        1031 => "0011001110110000",
        1032 => "0010110111010000",
        1033 => "0001111010100000",
        1034 => "0010100100000000",
        1035 => "0010101000000000",
        1036 => "0010010000110000",
        1037 => "0010100011110000",
        1038 => "0010011101010000",
        1039 => "0010100001100000",
        1040 => "0010111011100000",
        1041 => "0001110101100000",
        1042 => "0001101001110000",
        1043 => "0010110011100000",
        1044 => "0001111001010000",
        1045 => "0011011011000000",
        1046 => "0010011001100000",
        1047 => "0010000000110000",
        1048 => "0010010101110000",
        1049 => "0010011010100000",
        1050 => "0001111000110000",
        1051 => "0010100011100000",
        1052 => "0001111100010000",
        1053 => "0001100111100000",
        1054 => "0010101110000000",
        1055 => "0010101111110000",
        1056 => "0001101001110000",
        1057 => "0001111010100000",
        1058 => "0010111010010000",
        1059 => "0010011110110000",
        1060 => "0010111101110000",
        1061 => "0010110010100000",
        1062 => "0010110101110000",
        1063 => "0010100101000000",
        1064 => "0010101110100000",
        1065 => "0010001110100000",
        1066 => "0011000000110000",
        1067 => "0010100101010000",
        1068 => "0010100001010000",
        1069 => "0011000010010000",
        1070 => "0010111011010000",
        1071 => "0011011101010000",
        1072 => "0011110010000000",
        1073 => "0010110001100000",
        1074 => "0010101000000000",
        1075 => "0011100011000000",
        1076 => "0011000101010000",
        1077 => "0010100000000000",
        1078 => "0011100010110000",
        1079 => "0010011110110000",
        1080 => "0011000111110000",
        1081 => "0011001101000000",
        1082 => "0011010001010000",
        1083 => "0010111001100000",
        1084 => "0011100001100000",
        1085 => "0010101010010000",
        1086 => "0011100110000000",
        1087 => "0010111100100000",
        1088 => "0011001010000000",
        1089 => "0010100111000000",
        1090 => "0010010111100000",
        1091 => "0011011000010000",
        1092 => "0010110111110000",
        1093 => "0011010010100000",
        1094 => "0011010011100000",
        1095 => "0010110001100000",
        1096 => "0011000010110000",
        1097 => "0010110100010000",
        1098 => "0011100110010000",
        1099 => "0011010000010000",
        1100 => "0010110011010000",
        1101 => "0011010101110000",
        1102 => "0011000111110000",
        1103 => "0011000111110000",
        1104 => "0011010111000000",
        1105 => "0011101100100000",
        1106 => "0011001100010000",
        1107 => "0010111100000000",
        1108 => "0010100100110000",
        1109 => "0010001010100000",
        1110 => "0001111100000000",
        1111 => "0010001000110000",
        1112 => "0001111110100000",
        1113 => "0010000101110000",
        1114 => "0010000101110000",
        1115 => "0010000000110000",
        1116 => "0001010111110000",
        1117 => "0001110010000000",
        1118 => "0000001101000000",
        1119 => "0000110101100000",
        1120 => "0001011010100000",
        1121 => "0000011100000000",
        1122 => "0001000000110000",
        1123 => "0000110011010000",
        1124 => "0001000111010000",
        1125 => "0000101100100000",
        1126 => "0001100110010000",
        1127 => "0000111111000000",
        1128 => "0001011110010000",
        1129 => "0000111101100000",
        1130 => "0001110111000000",
        1131 => "0010010100100000",
        1132 => "0001101000000000",
        1133 => "0001011000000000",
        1134 => "0011001000110000",
        1135 => "0011000000000000",
        1136 => "0011000010110000",
        1137 => "0011100101010000",
        1138 => "0011101100110000",
        1139 => "0101000011100000",
        1140 => "0100101011110000",
        1141 => "0101111010010000",
        1142 => "0110100101110000",
        1143 => "0110101000110000",
        1144 => "0110000110010000",
        1145 => "0111000100110000",
        1146 => "1000101000010000",
        1147 => "0111011011010000",
        1148 => "1000001101110000",
        1149 => "1000101000100000",
        1150 => "1001000110000000",
        1151 => "1001110011110000",
        1152 => "1001100000000000",
        1153 => "1001000010000000",
        1154 => "1001101001110000",
        1155 => "1010001011100000",
        1156 => "1001110000100000",
        1157 => "1001111100000000",
        1158 => "1011000110110000",
        1159 => "1010010110000000",
        1160 => "1011000101010000",
        1161 => "1010100101000000",
        1162 => "1010101111100000",
        1163 => "1010110001110000",
        1164 => "1011010001100000",
        1165 => "1010110000000000",
        1166 => "1011111010000000",
        1167 => "1011100011110000",
        1168 => "1010101001110000",
        1169 => "1011101100010000",
        1170 => "1011010010100000",
        1171 => "1010111110000000",
        1172 => "1011100100110000",
        1173 => "1100001100100000",
        1174 => "1100001000010000",
        1175 => "1100001100000000",
        1176 => "1100011010100000",
        1177 => "1100011111000000",
        1178 => "1011110111110000",
        1179 => "1100100001110000",
        1180 => "1100101100000000",
        1181 => "1011111111100000",
        1182 => "1100000000110000",
        1183 => "1100001011000000",
        1184 => "1101011001110000",
        1185 => "1100010011110000",
        1186 => "1101100110100000",
        1187 => "1100010111010000",
        1188 => "1101011001010000",
        1189 => "1101001110100000",
        1190 => "1101000000000000",
        1191 => "1100110111000000",
        1192 => "1100011000000000",
        1193 => "1110011010110000",
        1194 => "1101011000010000",
        1195 => "1101110001010000",
        1196 => "1101111011000000",
        1197 => "1101011110100000",
        1198 => "1101100010000000",
        1199 => "1101000101110000",
        1200 => "1100110110100000",
        1201 => "1110000100010000",
        1202 => "1101010100110000",
        1203 => "1101010010100000",
        1204 => "1101001111100000",
        1205 => "1101000000110000",
        1206 => "1101011010110000",
        1207 => "1101011101100000",
        1208 => "1101101011010000",
        1209 => "1100111100010000",
        1210 => "1101111101010000",
        1211 => "1110010100000000",
        1212 => "1101011111010000",
        1213 => "1101101001100000",
        1214 => "1101001110010000",
        1215 => "1101110000010000",
        1216 => "1100110011000000",
        1217 => "1101110110110000",
        1218 => "1101011111100000",
        1219 => "1101101000010000",
        1220 => "1101101100010000",
        1221 => "1101111101000000",
        1222 => "1100011010010000",
        1223 => "1101011100010000",
        1224 => "1101110000010000",
        1225 => "1100100001100000",
        1226 => "1101000010100000",
        1227 => "1101010100110000",
        1228 => "1101100000000000",
        1229 => "1101000111010000",
        1230 => "1100011010000000",
        1231 => "1101100001000000",
        1232 => "1101001101000000",
        1233 => "1101011001010000",
        1234 => "1110001000010000",
        1235 => "1011110110010000",
        1236 => "1101000001010000",
        1237 => "1100100001000000",
        1238 => "1100111111100000",
        1239 => "1100100000000000",
        1240 => "1100110001100000",
        1241 => "1101001000110000",
        1242 => "1100101101100000",
        1243 => "1011111110010000",
        1244 => "1100110101110000",
        1245 => "1100011000010000",
        1246 => "1100101110100000",
        1247 => "1101000100010000",
        1248 => "1100101000100000",
        1249 => "1100101010010000",
        1250 => "1101100001100000",
        1251 => "1100111001110000",
        1252 => "1101011001000000",
        1253 => "1100011011110000",
        1254 => "1100010101010000",
        1255 => "1100100100000000",
        1256 => "1100101110010000",
        1257 => "1100010010010000",
        1258 => "1100111101000000",
        1259 => "1100111100110000",
        1260 => "1100011010110000",
        1261 => "1101001100100000",
        1262 => "1101010001110000",
        1263 => "1100111001110000",
        1264 => "1100111111100000",
        1265 => "1100010000000000",
        1266 => "1100111000010000",
        1267 => "1101100100010000",
        1268 => "1101001011110000",
        1269 => "1101100011100000",
        1270 => "1101100001000000",
        1271 => "1101111100110000",
        1272 => "1100110001100000",
        1273 => "1110101011000000",
        1274 => "1110000010010000",
        1275 => "1111000001100000",
        1276 => "1110101100110000",
        1277 => "1110100011010000",
        1278 => "1110111101010000",
        1279 => "1111000111110000",
        1280 => "1111001101010000",
        1281 => "1111100111010000",
        1282 => "1111111001100000",
        1283 => "1110111111100000",
        1284 => "1111000110110000",
        1285 => "1111100111000000",
        1286 => "1110011101110000",
        1287 => "1110111001000000",
        1288 => "1110101101010000",
        1289 => "1110011101110000",
        1290 => "1101111101010000",
        1291 => "1110101111000000",
        1292 => "1110001010000000",
        1293 => "1101100101010000",
        1294 => "1100100000100000",
        1295 => "1101001011110000",
        1296 => "1100010001100000",
        1297 => "1100000111010000",
        1298 => "1100000110100000",
        1299 => "1010111010000000",
        1300 => "1001100001110000",
        1301 => "1010000010010000",
        1302 => "1001111011110000",
        1303 => "1001000000000000",
        1304 => "1000100001000000",
        1305 => "1001100111000000",
        1306 => "0111101111110000",
        1307 => "1000100101010000",
        1308 => "0111000001100000",
        1309 => "0111011011000000",
        1310 => "0111100001010000",
        1311 => "0110110000100000",
        1312 => "0111000000100000",
        1313 => "0101111110010000",
        1314 => "0101100001100000",
        1315 => "0110000011100000",
        1316 => "0110000101110000",
        1317 => "0110001001010000",
        1318 => "0101100100110000",
        1319 => "0101001001100000",
        1320 => "0100101111010000",
        1321 => "0101010110010000",
        1322 => "0101000110010000",
        1323 => "0101110000100000",
        1324 => "0101010011100000",
        1325 => "0100111010100000",
        1326 => "0011111100110000",
        1327 => "0100010000000000",
        1328 => "0100101100000000",
        1329 => "0100111010000000",
        1330 => "0011101000110000",
        1331 => "0100001100010000",
        1332 => "0011010101100000",
        1333 => "0100010001000000",
        1334 => "0011111000000000",
        1335 => "0011101010010000",
        1336 => "0011110000110000",
        1337 => "0010111011000000",
        1338 => "0011011000110000",
        1339 => "0010111010010000",
        1340 => "0011000011100000",
        1341 => "0011101010110000",
        1342 => "0011010100110000",
        1343 => "0011000000100000",
        1344 => "0001110111100000",
        1345 => "0011011011100000",
        1346 => "0010010001000000",
        1347 => "0011011101000000",
        1348 => "0010010000110000",
        1349 => "0010011101110000",
        1350 => "0010011101010000",
        1351 => "0001110001000000",
        1352 => "0010110000010000",
        1353 => "0010110101010000",
        1354 => "0010110111000000",
        1355 => "0010100110110000",
        1356 => "0010000101110000",
        1357 => "0001101011000000",
        1358 => "0011001100110000",
        1359 => "0010010001010000",
        1360 => "0010111001000000",
        1361 => "0001111101110000",
        1362 => "0010001011000000",
        1363 => "0011000111000000",
        1364 => "0010001001000000",
        1365 => "0001110001110000",
        1366 => "0010101101110000",
        1367 => "0001111010000000",
        1368 => "0010000001100000",
        1369 => "0011001000100000",
        1370 => "0011001110100000",
        1371 => "0001110101010000",
        1372 => "0010100111100000",
        1373 => "0010101100100000",
        1374 => "0010100110110000",
        1375 => "0010011100110000",
        1376 => "0010000110000000",
        1377 => "0001101110000000",
        1378 => "0010010111010000",
        1379 => "0010101000010000",
        1380 => "0010101010100000",
        1381 => "0011000000010000",
        1382 => "0010011100000000",
        1383 => "0011000010110000",
        1384 => "0010011010000000",
        1385 => "0010001100110000",
        1386 => "0010100000000000",
        1387 => "0010101100110000",
        1388 => "0010010000000000",
        1389 => "0010011110010000",
        1390 => "0011000010110000",
        1391 => "0011100001110000",
        1392 => "0010100011010000",
        1393 => "0010100111010000",
        1394 => "0010111000000000",
        1395 => "0010110111000000",
        1396 => "0011010001100000",
        1397 => "0011010001100000",
        1398 => "0010001110000000",
        1399 => "0011001010000000",
        1400 => "0010100001000000",
        1401 => "0010110100110000",
        1402 => "0010111011000000",
        1403 => "0011011110100000",
        1404 => "0011001001010000",
        1405 => "0010000001000000",
        1406 => "0010111111110000",
        1407 => "0010111010100000",
        1408 => "0011001000010000",
        1409 => "0010011110100000",
        1410 => "0010101010000000",
        1411 => "0010111000110000",
        1412 => "0011000100000000",
        1413 => "0011100100110000",
        1414 => "0011010000000000",
        1415 => "0011000101110000",
        1416 => "0011110011110000",
        1417 => "0010111100100000",
        1418 => "0010110101110000",
        1419 => "0010101010100000",
        1420 => "0010110000010000",
        1421 => "0011000110000000",
        1422 => "0011101001100000",
        1423 => "0011000010100000",
        1424 => "0011010010100000",
        1425 => "0011010010010000",
        1426 => "0010111010000000",
        1427 => "0010101100010000",
        1428 => "0011000100100000",
        1429 => "0001111010100000",
        1430 => "0010010000110000",
        1431 => "0001111101110000",
        1432 => "0010011111110000",
        1433 => "0001111111110000",
        1434 => "0001010100110000",
        1435 => "0001010011100000",
        1436 => "0001110111110000",
        1437 => "0001000000010000",
        1438 => "0001000100110000",
        1439 => "0000101110100000",
        1440 => "0000101101110000",
        1441 => "0000100011010000",
        1442 => "0001010011100000",
        1443 => "0000101111100000",
        1444 => "0000000000000000",
        1445 => "0001000010100000",
        1446 => "0000101010110000",
        1447 => "0001001110110000",
        1448 => "0000010011010000",
        1449 => "0010000110110000",
        1450 => "0001000001000000",
        1451 => "0001110111110000",
        1452 => "0001000100110000",
        1453 => "0001111110000000",
        1454 => "0011000110110000",
        1455 => "0010111111000000",
        1456 => "0011000100100000",
        1457 => "0011100000010000",
        1458 => "0100110100000000",
        1459 => "0011101111010000",
        1460 => "0101010100000000",
        1461 => "0101010101110000",
        1462 => "0110000100100000",
        1463 => "0110011101010000",
        1464 => "0110111001100000",
        1465 => "0110110001110000",
        1466 => "1000001011010000",
        1467 => "1000100011100000",
        1468 => "0111111101000000",
        1469 => "1000110101100000",
        1470 => "1000101110110000",
        1471 => "1000101011010000",
        1472 => "1010000110010000",
        1473 => "1001010101000000",
        1474 => "1010001001000000",
        1475 => "1001100001110000",
        1476 => "1010000111110000",
        1477 => "1001101110110000",
        1478 => "1010110001110000",
        1479 => "1010011110010000",
        1480 => "1010011010110000",
        1481 => "1100011111010000",
        1482 => "1011011110010000",
        1483 => "1011110011100000",
        1484 => "1010111101100000",
        1485 => "1010111101100000",
        1486 => "1010110100110000",
        1487 => "1011010101010000",
        1488 => "1011001100100000",
        1489 => "1011110000110000",
        1490 => "1100011001100000",
        1491 => "1011101111000000",
        1492 => "1100011010110000",
        1493 => "1100001010010000",
        1494 => "1100110111100000",
        1495 => "1011110000010000",
        1496 => "1011110110000000",
        1497 => "1011101111100000",
        1498 => "1100000011000000",
        1499 => "1100011100000000",
        1500 => "1100110011000000",
        1501 => "1101000011110000",
        1502 => "1101000010000000",
        1503 => "1101001111100000",
        1504 => "1100111011110000",
        1505 => "1101001100100000",
        1506 => "1100001100000000",
        1507 => "1101001001100000",
        1508 => "1101011011100000",
        1509 => "1101001001010000",
        1510 => "1101101011010000",
        1511 => "1101001111100000",
        1512 => "1100110111000000",
        1513 => "1101010101010000",
        1514 => "1101010110110000",
        1515 => "1101010011010000",
        1516 => "1101001111100000",
        1517 => "1101111001110000",
        1518 => "1100100100110000",
        1519 => "1101101001000000",
        1520 => "1101001010000000",
        1521 => "1101101000010000",
        1522 => "1110000101110000",
        1523 => "1110001011100000",
        1524 => "1101100000010000",
        1525 => "1101100001100000",
        1526 => "1101111110100000",
        1527 => "1101110111000000",
        1528 => "1101100100110000",
        1529 => "1101001110100000",
        1530 => "1101011101010000",
        1531 => "1110000111010000",
        1532 => "1100110100110000",
        1533 => "1101100001100000",
        1534 => "1101000101100000",
        1535 => "1101111111000000",
        1536 => "1101010101100000",
        1537 => "1101100011110000",
        1538 => "1100110101000000",
        1539 => "1101100111100000",
        1540 => "1101010011000000",
        1541 => "1101100100000000",
        1542 => "1101110001100000",
        1543 => "1101000101100000",
        1544 => "1101100111000000",
        1545 => "1101001011000000",
        1546 => "1100100101110000",
        1547 => "1100110111000000",
        1548 => "1101001011100000",
        1549 => "1101011001000000",
        1550 => "1101100111110000",
        1551 => "1110000001110000",
        1552 => "1100111000100000",
        1553 => "1101000001100000",
        1554 => "1101001100000000",
        1555 => "1100011010110000",
        1556 => "1100001110110000",
        1557 => "1100100110100000",
        1558 => "1100101011110000",
        1559 => "1100110101110000",
        1560 => "1101010111110000",
        1561 => "1101001100100000",
        1562 => "1100111001010000",
        1563 => "1100010110100000",
        1564 => "1100010011000000",
        1565 => "1101010001010000",
        1566 => "1101011001100000",
        1567 => "1011111010100000",
        1568 => "1100100101100000",
        1569 => "1100011111100000",
        1570 => "1101100000100000",
        1571 => "1100111011000000",
        1572 => "1011100100100000",
        1573 => "1100011001100000",
        1574 => "1101001000110000",
        1575 => "1101000000100000",
        1576 => "1100010000000000",
        1577 => "1100100110000000",
        1578 => "1101000000000000",
        1579 => "1100001011010000",
        1580 => "1100101100100000",
        1581 => "1100011110010000",
        1582 => "1100001010010000",
        1583 => "1100101100000000",
        1584 => "1101001100100000",
        1585 => "1100000101100000",
        1586 => "1100011010010000",
        1587 => "1101011011010000",
        1588 => "1101000110100000",
        1589 => "1101010101000000",
        1590 => "1101011111100000",
        1591 => "1110010001000000",
        1592 => "1110010110010000",
        1593 => "1101100111110000",
        1594 => "1110001100110000",
        1595 => "1110110110000000",
        1596 => "1110010001110000",
        1597 => "1101101100000000",
        1598 => "1110111100000000",
        1599 => "1110111011000000"
    );
BEGIN
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            data_out <= rom(address);
        END IF;
    END PROCESS;
END Behavioral;