-- megafunction wizard: %RAM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: data_mem.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.0 Build 208 07/03/2011 SP 1 SJ Full Version
-- ************************************************************
--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.

-- Zoran Salcic

library ieee;
use ieee.std_logic_1164.all;

library altera_mf;
use altera_mf.all;

entity data_mem is
	port (
		address : in std_logic_vector (13 downto 0);
		clock   : in std_logic := '1';
		data    : in std_logic_vector (15 downto 0);
		wren    : in std_logic;
		q       : out std_logic_vector (15 downto 0)
	);
end data_mem;
architecture SYN of data_mem is

	signal sub_wire0 : std_logic_vector (15 downto 0);

	component altsyncram
		generic (
			clock_enable_input_a   : string;
			clock_enable_output_a  : string;
			intended_device_family : string;
			lpm_hint               : string;
			lpm_type               : string;
			numwords_a             : natural;
			operation_mode         : string;
			outdata_aclr_a         : string;
			outdata_reg_a          : string;
			power_up_uninitialized : string;
			ram_block_type         : string;
			widthad_a              : natural;
			width_a                : natural;
			width_byteena_a        : natural
		);
		port (
			address_a : in std_logic_vector (13 downto 0);
			clock0    : in std_logic;
			data_a    : in std_logic_vector (15 downto 0);
			wren_a    : in std_logic;
			q_a       : out std_logic_vector (15 downto 0)
		);
	end component;

begin
	q <= sub_wire0(15 downto 0);

	altsyncram_component : altsyncram
	generic map(
		clock_enable_input_a   => "BYPASS",
		clock_enable_output_a  => "BYPASS",
		intended_device_family => "Cyclone II",
		lpm_hint               => "ENABLE_RUNTIME_MOD=NO",
		lpm_type               => "altsyncram",
		numwords_a             => 4096,
		operation_mode         => "SINGLE_PORT",
		outdata_aclr_a         => "NONE",
		outdata_reg_a          => "UNREGISTERED",
		power_up_uninitialized => "FALSE",
		ram_block_type         => "M4K",
		widthad_a              => 14,
		width_a                => 16,
		width_byteena_a        => 1
	)
	port map(
		clock0    => clock,
		address_a => address,
		data_a    => data,
		wren_a    => wren,
		q_a       => sub_wire0
	);

end SYN;