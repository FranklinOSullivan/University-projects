LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY wave IS
    PORT (
        clk : IN STD_LOGIC;
        address : IN INTEGER RANGE 0 TO 1599; -- 10 cycles * 16000 samples/s / 50 Hz
        data_out : OUT unsigned(15 DOWNTO 0) -- 8-bit output
    );
END wave;

ARCHITECTURE beh OF wave IS
    TYPE rom_type IS ARRAY (0 TO 1599) OF unsigned(15 DOWNTO 0);
    ---FAT array with 1600 samples of the power signal
    SIGNAL rom : rom_type := (
         0 => "1100110010010000",
    1 => "1100101010000000",
    2 => "1100100010000000",
    3 => "1100011001100000",
    4 => "1100010001000000",
    5 => "1100001000100000",
    6 => "1100000000000000",
    7 => "1011110111010000",
    8 => "1011101110010000",
    9 => "1011100101010000",
    10 => "1011011100010000",
    11 => "1011010011010000",
    12 => "1011001010000000",
    13 => "1011000000110000",
    14 => "1010110111100000",
    15 => "1010101110000000",
    16 => "1010100100100000",
    17 => "1010011011000000",
    18 => "1010010001010000",
    19 => "1010000111110000",
    20 => "1001111110000000",
    21 => "1001110100010000",
    22 => "1001101010100000",
    23 => "1001100000100000",
    24 => "1001010110110000",
    25 => "1001001100110000",
    26 => "1001000010110000",
    27 => "1000111000110000",
    28 => "1000101110110000",
    29 => "1000100100110000",
    30 => "1000011010110000",
    31 => "1000010000110000",
    32 => "1000000110110000",
    33 => "0111111100100000",
    34 => "0111110010100000",
    35 => "0111101000100000",
    36 => "0111011110100000",
    37 => "0111010100100000",
    38 => "0111001010100000",
    39 => "0111000000100000",
    40 => "0110110110100000",
    41 => "0110101100100000",
    42 => "0110100010110000",
    43 => "0110011000110000",
    44 => "0110001111000000",
    45 => "0110000101010000",
    46 => "0101111011100000",
    47 => "0101110001110000",
    48 => "0101101000010000",
    49 => "0101011110100000",
    50 => "0101010101000000",
    51 => "0101001011110000",
    52 => "0101000010010000",
    53 => "0100111001000000",
    54 => "0100101111110000",
    55 => "0100100110100000",
    56 => "0100011101100000",
    57 => "0100010100100000",
    58 => "0100001011110000",
    59 => "0100000011000000",
    60 => "0011111010010000",
    61 => "0011110001110000",
    62 => "0011101001010000",
    63 => "0011100000110000",
    64 => "0011011000100000",
    65 => "0011010000010000",
    66 => "0011001000010000",
    67 => "0011000000100000",
    68 => "0010111000110000",
    69 => "0010110001000000",
    70 => "0010101001100000",
    71 => "0010100010000000",
    72 => "0010011010110000",
    73 => "0010010011100000",
    74 => "0010001100110000",
    75 => "0010000101110000",
    76 => "0001111111000000",
    77 => "0001111000100000",
    78 => "0001110010000000",
    79 => "0001101100000000",
    80 => "0001100101110000",
    81 => "0001011111110000",
    82 => "0001011010000000",
    83 => "0001010100100000",
    84 => "0001001111000000",
    85 => "0001001001110000",
    86 => "0001000100100000",
    87 => "0000111111110000",
    88 => "0000111011000000",
    89 => "0000110110010000",
    90 => "0000110010000000",
    91 => "0000101101110000",
    92 => "0000101001100000",
    93 => "0000100101110000",
    94 => "0000100010000000",
    95 => "0000011110100000",
    96 => "0000011011010000",
    97 => "0000011000000000",
    98 => "0000010101000000",
    99 => "0000010010010000",
    100 => "0000001111110000",
    101 => "0000001101100000",
    102 => "0000001011010000",
    103 => "0000001001010000",
    104 => "0000000111100000",
    105 => "0000000101110000",
    106 => "0000000100100000",
    107 => "0000000011010000",
    108 => "0000000010010000",
    109 => "0000000001010000",
    110 => "0000000000110000",
    111 => "0000000000010000",
    112 => "0000000000000000",
    113 => "0000000000000000",
    114 => "0000000000010000",
    115 => "0000000000100000",
    116 => "0000000001000000",
    117 => "0000000001110000",
    118 => "0000000010110000",
    119 => "0000000100000000",
    120 => "0000000101010000",
    121 => "0000000110110000",
    122 => "0000001000100000",
    123 => "0000001010100000",
    124 => "0000001100100000",
    125 => "0000001111000000",
    126 => "0000010001100000",
    127 => "0000010100000000",
    128 => "0000010111000000",
    129 => "0000011010000000",
    130 => "0000011101010000",
    131 => "0000100000110000",
    132 => "0000100100100000",
    133 => "0000101000010000",
    134 => "0000101100010000",
    135 => "0000110000100000",
    136 => "0000110100110000",
    137 => "0000111001010000",
    138 => "0000111110000000",
    139 => "0001000010110000",
    140 => "0001001000000000",
    141 => "0001001101010000",
    142 => "0001010010100000",
    143 => "0001011000000000",
    144 => "0001011101110000",
    145 => "0001100011110000",
    146 => "0001101001110000",
    147 => "0001110000000000",
    148 => "0001110110010000",
    149 => "0001111100110000",
    150 => "0010000011100000",
    151 => "0010001010010000",
    152 => "0010010001010000",
    153 => "0010011000010000",
    154 => "0010011111100000",
    155 => "0010100110110000",
    156 => "0010101110010000",
    157 => "0010110110000000",
    158 => "0010111101110000",
    159 => "0011000101100000",
    160 => "0011001101100000",
    161 => "0011010101110000",
    162 => "0011011101110000",
    163 => "0011100110010000",
    164 => "0011101110110000",
    165 => "0011110111010000",
    166 => "0011111111110000",
    167 => "0100001000100000",
    168 => "0100010001100000",
    169 => "0100011010100000",
    170 => "0100100011100000",
    171 => "0100101100100000",
    172 => "0100110101110000",
    173 => "0100111111000000",
    174 => "0101001000010000",
    175 => "0101010001110000",
    176 => "0101011011010000",
    177 => "0101100100110000",
    178 => "0101101110100000",
    179 => "0101111000000000",
    180 => "0110000001110000",
    181 => "0110001011100000",
    182 => "0110010101010000",
    183 => "0110011111010000",
    184 => "0110101001000000",
    185 => "0110110011000000",
    186 => "0110111101000000",
    187 => "0111000111000000",
    188 => "0111010001000000",
    189 => "0111011011000000",
    190 => "0111100101000000",
    191 => "0111101111000000",
    192 => "0111111001000000",
    193 => "1000000011010000",
    194 => "1000001101010000",
    195 => "1000010111010000",
    196 => "1000100001010000",
    197 => "1000101011010000",
    198 => "1000110101010000",
    199 => "1000111111010000",
    200 => "1001001001010000",
    201 => "1001010011010000",
    202 => "1001011101000000",
    203 => "1001100111000000",
    204 => "1001110000110000",
    205 => "1001111010100000",
    206 => "1010000100010000",
    207 => "1010001110000000",
    208 => "1010010111100000",
    209 => "1010100001010000",
    210 => "1010101010110000",
    211 => "1010110100000000",
    212 => "1010111101100000",
    213 => "1011000110110000",
    214 => "1011010000000000",
    215 => "1011011001010000",
    216 => "1011100010010000",
    217 => "1011101011010000",
    218 => "1011110100000000",
    219 => "1011111100110000",
    220 => "1100000101100000",
    221 => "1100001110000000",
    222 => "1100010110100000",
    223 => "1100011111000000",
    224 => "1100100111010000",
    225 => "1100101111100000",
    226 => "1100110111100000",
    227 => "1100111111010000",
    228 => "1101000111000000",
    229 => "1101001110110000",
    230 => "1101010110010000",
    231 => "1101011101110000",
    232 => "1101100101000000",
    233 => "1101101100010000",
    234 => "1101110011000000",
    235 => "1101111010000000",
    236 => "1110000000110000",
    237 => "1110000111010000",
    238 => "1110001101110000",
    239 => "1110010011110000",
    240 => "1110011010000000",
    241 => "1110100000000000",
    242 => "1110100101110000",
    243 => "1110101011010000",
    244 => "1110110000110000",
    245 => "1110110110000000",
    246 => "1110111011010000",
    247 => "1111000000000000",
    248 => "1111000100110000",
    249 => "1111001001100000",
    250 => "1111001101110000",
    251 => "1111010010000000",
    252 => "1111010110010000",
    253 => "1111011010000000",
    254 => "1111011101110000",
    255 => "1111100001010000",
    256 => "1111100100100000",
    257 => "1111100111110000",
    258 => "1111101010110000",
    259 => "1111101101100000",
    260 => "1111110000000000",
    261 => "1111110010010000",
    262 => "1111110100100000",
    263 => "1111110110100000",
    264 => "1111111000010000",
    265 => "1111111010000000",
    266 => "1111111011010000",
    267 => "1111111100100000",
    268 => "1111111101100000",
    269 => "1111111110100000",
    270 => "1111111111000000",
    271 => "1111111111100000",
    272 => "1111111111110000",
    273 => "1111111111110000",
    274 => "1111111111100000",
    275 => "1111111111010000",
    276 => "1111111110110000",
    277 => "1111111110000000",
    278 => "1111111101000000",
    279 => "1111111011110000",
    280 => "1111111010100000",
    281 => "1111111001000000",
    282 => "1111110111010000",
    283 => "1111110101010000",
    284 => "1111110011010000",
    285 => "1111110000110000",
    286 => "1111101110010000",
    287 => "1111101011110000",
    288 => "1111101000110000",
    289 => "1111100101110000",
    290 => "1111100010100000",
    291 => "1111011111000000",
    292 => "1111011011010000",
    293 => "1111010111100000",
    294 => "1111010011100000",
    295 => "1111001111010000",
    296 => "1111001011000000",
    297 => "1111000110100000",
    298 => "1111000001110000",
    299 => "1110111101000000",
    300 => "1110110111110000",
    301 => "1110110010100000",
    302 => "1110101101010000",
    303 => "1110100111110000",
    304 => "1110100010000000",
    305 => "1110011100000000",
    306 => "1110010110000000",
    307 => "1110001111110000",
    308 => "1110001001100000",
    309 => "1110000011000000",
    310 => "1101111100010000",
    311 => "1101110101100000",
    312 => "1101101110100000",
    313 => "1101100111100000",
    314 => "1101100000010000",
    315 => "1101011001000000",
    316 => "1101010001100000",
    317 => "1101001001110000",
    318 => "1101000010000000",
    319 => "1100111010010000",
    320 => "1100110010010000",
    321 => "1100101010000000",
    322 => "1100100010000000",
    323 => "1100011001100000",
    324 => "1100010001000000",
    325 => "1100001000100000",
    326 => "1100000000000000",
    327 => "1011110111010000",
    328 => "1011101110010000",
    329 => "1011100101010000",
    330 => "1011011100010000",
    331 => "1011010011010000",
    332 => "1011001010000000",
    333 => "1011000000110000",
    334 => "1010110111100000",
    335 => "1010101110000000",
    336 => "1010100100100000",
    337 => "1010011011000000",
    338 => "1010010001010000",
    339 => "1010000111110000",
    340 => "1001111110000000",
    341 => "1001110100010000",
    342 => "1001101010100000",
    343 => "1001100000100000",
    344 => "1001010110110000",
    345 => "1001001100110000",
    346 => "1001000010110000",
    347 => "1000111000110000",
    348 => "1000101110110000",
    349 => "1000100100110000",
    350 => "1000011010110000",
    351 => "1000010000110000",
    352 => "1000000110110000",
    353 => "0111111100100000",
    354 => "0111110010100000",
    355 => "0111101000100000",
    356 => "0111011110100000",
    357 => "0111010100100000",
    358 => "0111001010100000",
    359 => "0111000000100000",
    360 => "0110110110100000",
    361 => "0110101100100000",
    362 => "0110100010110000",
    363 => "0110011000110000",
    364 => "0110001111000000",
    365 => "0110000101010000",
    366 => "0101111011100000",
    367 => "0101110001110000",
    368 => "0101101000010000",
    369 => "0101011110100000",
    370 => "0101010101000000",
    371 => "0101001011110000",
    372 => "0101000010010000",
    373 => "0100111001000000",
    374 => "0100101111110000",
    375 => "0100100110100000",
    376 => "0100011101100000",
    377 => "0100010100100000",
    378 => "0100001011110000",
    379 => "0100000011000000",
    380 => "0011111010010000",
    381 => "0011110001110000",
    382 => "0011101001010000",
    383 => "0011100000110000",
    384 => "0011011000100000",
    385 => "0011010000010000",
    386 => "0011001000010000",
    387 => "0011000000100000",
    388 => "0010111000110000",
    389 => "0010110001000000",
    390 => "0010101001100000",
    391 => "0010100010000000",
    392 => "0010011010110000",
    393 => "0010010011100000",
    394 => "0010001100110000",
    395 => "0010000101110000",
    396 => "0001111111000000",
    397 => "0001111000100000",
    398 => "0001110010000000",
    399 => "0001101100000000",
    400 => "0001100101110000",
    401 => "0001011111110000",
    402 => "0001011010000000",
    403 => "0001010100100000",
    404 => "0001001111000000",
    405 => "0001001001110000",
    406 => "0001000100100000",
    407 => "0000111111110000",
    408 => "0000111011000000",
    409 => "0000110110010000",
    410 => "0000110010000000",
    411 => "0000101101110000",
    412 => "0000101001100000",
    413 => "0000100101110000",
    414 => "0000100010000000",
    415 => "0000011110100000",
    416 => "0000011011010000",
    417 => "0000011000000000",
    418 => "0000010101000000",
    419 => "0000010010010000",
    420 => "0000001111110000",
    421 => "0000001101100000",
    422 => "0000001011010000",
    423 => "0000001001010000",
    424 => "0000000111100000",
    425 => "0000000101110000",
    426 => "0000000100100000",
    427 => "0000000011010000",
    428 => "0000000010010000",
    429 => "0000000001010000",
    430 => "0000000000110000",
    431 => "0000000000010000",
    432 => "0000000000000000",
    433 => "0000000000000000",
    434 => "0000000000010000",
    435 => "0000000000100000",
    436 => "0000000001000000",
    437 => "0000000001110000",
    438 => "0000000010110000",
    439 => "0000000100000000",
    440 => "0000000101010000",
    441 => "0000000110110000",
    442 => "0000001000100000",
    443 => "0000001010100000",
    444 => "0000001100100000",
    445 => "0000001111000000",
    446 => "0000010001100000",
    447 => "0000010100000000",
    448 => "0000010111000000",
    449 => "0000011010000000",
    450 => "0000011101010000",
    451 => "0000100000110000",
    452 => "0000100100100000",
    453 => "0000101000010000",
    454 => "0000101100010000",
    455 => "0000110000100000",
    456 => "0000110100110000",
    457 => "0000111001010000",
    458 => "0000111110000000",
    459 => "0001000010110000",
    460 => "0001001000000000",
    461 => "0001001101010000",
    462 => "0001010010100000",
    463 => "0001011000000000",
    464 => "0001011101110000",
    465 => "0001100011110000",
    466 => "0001101001110000",
    467 => "0001110000000000",
    468 => "0001110110010000",
    469 => "0001111100110000",
    470 => "0010000011100000",
    471 => "0010001010010000",
    472 => "0010010001010000",
    473 => "0010011000010000",
    474 => "0010011111100000",
    475 => "0010100110110000",
    476 => "0010101110010000",
    477 => "0010110110000000",
    478 => "0010111101110000",
    479 => "0011000101100000",
    480 => "0011001101100000",
    481 => "0011010101110000",
    482 => "0011011101110000",
    483 => "0011100110010000",
    484 => "0011101110110000",
    485 => "0011110111010000",
    486 => "0011111111110000",
    487 => "0100001000100000",
    488 => "0100010001100000",
    489 => "0100011010100000",
    490 => "0100100011100000",
    491 => "0100101100100000",
    492 => "0100110101110000",
    493 => "0100111111000000",
    494 => "0101001000010000",
    495 => "0101010001110000",
    496 => "0101011011010000",
    497 => "0101100100110000",
    498 => "0101101110100000",
    499 => "0101111000000000",
    500 => "0110000001110000",
    501 => "0110001011100000",
    502 => "0110010101010000",
    503 => "0110011111010000",
    504 => "0110101001000000",
    505 => "0110110011000000",
    506 => "0110111101000000",
    507 => "0111000111000000",
    508 => "0111010001000000",
    509 => "0111011011000000",
    510 => "0111100101000000",
    511 => "0111101111000000",
    512 => "0111111001000000",
    513 => "1000000011010000",
    514 => "1000001101010000",
    515 => "1000010111010000",
    516 => "1000100001010000",
    517 => "1000101011010000",
    518 => "1000110101010000",
    519 => "1000111111010000",
    520 => "1001001001010000",
    521 => "1001010011010000",
    522 => "1001011101000000",
    523 => "1001100111000000",
    524 => "1001110000110000",
    525 => "1001111010100000",
    526 => "1010000100010000",
    527 => "1010001110000000",
    528 => "1010010111100000",
    529 => "1010100001010000",
    530 => "1010101010110000",
    531 => "1010110100000000",
    532 => "1010111101100000",
    533 => "1011000110110000",
    534 => "1011010000000000",
    535 => "1011011001010000",
    536 => "1011100010010000",
    537 => "1011101011010000",
    538 => "1011110100000000",
    539 => "1011111100110000",
    540 => "1100000101100000",
    541 => "1100001110000000",
    542 => "1100010110100000",
    543 => "1100011111000000",
    544 => "1100100111010000",
    545 => "1100101111100000",
    546 => "1100110111100000",
    547 => "1100111111010000",
    548 => "1101000111000000",
    549 => "1101001110110000",
    550 => "1101010110010000",
    551 => "1101011101110000",
    552 => "1101100101000000",
    553 => "1101101100010000",
    554 => "1101110011000000",
    555 => "1101111010000000",
    556 => "1110000000110000",
    557 => "1110000111010000",
    558 => "1110001101110000",
    559 => "1110010011110000",
    560 => "1110011010000000",
    561 => "1110100000000000",
    562 => "1110100101110000",
    563 => "1110101011010000",
    564 => "1110110000110000",
    565 => "1110110110000000",
    566 => "1110111011010000",
    567 => "1111000000000000",
    568 => "1111000100110000",
    569 => "1111001001100000",
    570 => "1111001101110000",
    571 => "1111010010000000",
    572 => "1111010110010000",
    573 => "1111011010000000",
    574 => "1111011101110000",
    575 => "1111100001010000",
    576 => "1111100100100000",
    577 => "1111100111110000",
    578 => "1111101010110000",
    579 => "1111101101100000",
    580 => "1111110000000000",
    581 => "1111110010010000",
    582 => "1111110100100000",
    583 => "1111110110100000",
    584 => "1111111000010000",
    585 => "1111111010000000",
    586 => "1111111011010000",
    587 => "1111111100100000",
    588 => "1111111101100000",
    589 => "1111111110100000",
    590 => "1111111111000000",
    591 => "1111111111100000",
    592 => "1111111111110000",
    593 => "1111111111110000",
    594 => "1111111111100000",
    595 => "1111111111010000",
    596 => "1111111110110000",
    597 => "1111111110000000",
    598 => "1111111101000000",
    599 => "1111111011110000",
    600 => "1111111010100000",
    601 => "1111111001000000",
    602 => "1111110111010000",
    603 => "1111110101010000",
    604 => "1111110011010000",
    605 => "1111110000110000",
    606 => "1111101110010000",
    607 => "1111101011110000",
    608 => "1111101000110000",
    609 => "1111100101110000",
    610 => "1111100010100000",
    611 => "1111011111000000",
    612 => "1111011011010000",
    613 => "1111010111100000",
    614 => "1111010011100000",
    615 => "1111001111010000",
    616 => "1111001011000000",
    617 => "1111000110100000",
    618 => "1111000001110000",
    619 => "1110111101000000",
    620 => "1110110111110000",
    621 => "1110110010100000",
    622 => "1110101101010000",
    623 => "1110100111110000",
    624 => "1110100010000000",
    625 => "1110011100000000",
    626 => "1110010110000000",
    627 => "1110001111110000",
    628 => "1110001001100000",
    629 => "1110000011000000",
    630 => "1101111100010000",
    631 => "1101110101100000",
    632 => "1101101110100000",
    633 => "1101100111100000",
    634 => "1101100000010000",
    635 => "1101011001000000",
    636 => "1101010001100000",
    637 => "1101001001110000",
    638 => "1101000010000000",
    639 => "1100111010010000",
    640 => "1100110010010000",
    641 => "1100101010000000",
    642 => "1100100010000000",
    643 => "1100011001100000",
    644 => "1100010001000000",
    645 => "1100001000100000",
    646 => "1100000000000000",
    647 => "1011110111010000",
    648 => "1011101110010000",
    649 => "1011100101010000",
    650 => "1011011100010000",
    651 => "1011010011010000",
    652 => "1011001010000000",
    653 => "1011000000110000",
    654 => "1010110111100000",
    655 => "1010101110000000",
    656 => "1010100100100000",
    657 => "1010011011000000",
    658 => "1010010001010000",
    659 => "1010000111110000",
    660 => "1001111110000000",
    661 => "1001110100010000",
    662 => "1001101010100000",
    663 => "1001100000100000",
    664 => "1001010110110000",
    665 => "1001001100110000",
    666 => "1001000010110000",
    667 => "1000111000110000",
    668 => "1000101110110000",
    669 => "1000100100110000",
    670 => "1000011010110000",
    671 => "1000010000110000",
    672 => "1000000110110000",
    673 => "0111111100100000",
    674 => "0111110010100000",
    675 => "0111101000100000",
    676 => "0111011110100000",
    677 => "0111010100100000",
    678 => "0111001010100000",
    679 => "0111000000100000",
    680 => "0110110110100000",
    681 => "0110101100100000",
    682 => "0110100010110000",
    683 => "0110011000110000",
    684 => "0110001111000000",
    685 => "0110000101010000",
    686 => "0101111011100000",
    687 => "0101110001110000",
    688 => "0101101000010000",
    689 => "0101011110100000",
    690 => "0101010101000000",
    691 => "0101001011110000",
    692 => "0101000010010000",
    693 => "0100111001000000",
    694 => "0100101111110000",
    695 => "0100100110100000",
    696 => "0100011101100000",
    697 => "0100010100100000",
    698 => "0100001011110000",
    699 => "0100000011000000",
    700 => "0011111010010000",
    701 => "0011110001110000",
    702 => "0011101001010000",
    703 => "0011100000110000",
    704 => "0011011000100000",
    705 => "0011010000010000",
    706 => "0011001000010000",
    707 => "0011000000100000",
    708 => "0010111000110000",
    709 => "0010110001000000",
    710 => "0010101001100000",
    711 => "0010100010000000",
    712 => "0010011010110000",
    713 => "0010010011100000",
    714 => "0010001100110000",
    715 => "0010000101110000",
    716 => "0001111111000000",
    717 => "0001111000100000",
    718 => "0001110010000000",
    719 => "0001101100000000",
    720 => "0001100101110000",
    721 => "0001011111110000",
    722 => "0001011010000000",
    723 => "0001010100100000",
    724 => "0001001111000000",
    725 => "0001001001110000",
    726 => "0001000100100000",
    727 => "0000111111110000",
    728 => "0000111011000000",
    729 => "0000110110010000",
    730 => "0000110010000000",
    731 => "0000101101110000",
    732 => "0000101001100000",
    733 => "0000100101110000",
    734 => "0000100010000000",
    735 => "0000011110100000",
    736 => "0000011011010000",
    737 => "0000011000000000",
    738 => "0000010101000000",
    739 => "0000010010010000",
    740 => "0000001111110000",
    741 => "0000001101100000",
    742 => "0000001011010000",
    743 => "0000001001010000",
    744 => "0000000111100000",
    745 => "0000000101110000",
    746 => "0000000100100000",
    747 => "0000000011010000",
    748 => "0000000010010000",
    749 => "0000000001010000",
    750 => "0000000000110000",
    751 => "0000000000010000",
    752 => "0000000000000000",
    753 => "0000000000000000",
    754 => "0000000000010000",
    755 => "0000000000100000",
    756 => "0000000001000000",
    757 => "0000000001110000",
    758 => "0000000010110000",
    759 => "0000000100000000",
    760 => "0000000101010000",
    761 => "0000000110110000",
    762 => "0000001000100000",
    763 => "0000001010100000",
    764 => "0000001100100000",
    765 => "0000001111000000",
    766 => "0000010001100000",
    767 => "0000010100000000",
    768 => "0000010111000000",
    769 => "0000011010000000",
    770 => "0000011101010000",
    771 => "0000100000110000",
    772 => "0000100100100000",
    773 => "0000101000010000",
    774 => "0000101100010000",
    775 => "0000110000100000",
    776 => "0000110100110000",
    777 => "0000111001010000",
    778 => "0000111110000000",
    779 => "0001000010110000",
    780 => "0001001000000000",
    781 => "0001001101010000",
    782 => "0001010010100000",
    783 => "0001011000000000",
    784 => "0001011101110000",
    785 => "0001100011110000",
    786 => "0001101001110000",
    787 => "0001110000000000",
    788 => "0001110110010000",
    789 => "0001111100110000",
    790 => "0010000011100000",
    791 => "0010001010010000",
    792 => "0010010001010000",
    793 => "0010011000010000",
    794 => "0010011111100000",
    795 => "0010100110110000",
    796 => "0010101110010000",
    797 => "0010110110000000",
    798 => "0010111101110000",
    799 => "0011000101100000",
    800 => "0011001101100000",
    801 => "0011010101110000",
    802 => "0011011101110000",
    803 => "0011100110010000",
    804 => "0011101110110000",
    805 => "0011110111010000",
    806 => "0011111111110000",
    807 => "0100001000100000",
    808 => "0100010001100000",
    809 => "0100011010100000",
    810 => "0100100011100000",
    811 => "0100101100100000",
    812 => "0100110101110000",
    813 => "0100111111000000",
    814 => "0101001000010000",
    815 => "0101010001110000",
    816 => "0101011011010000",
    817 => "0101100100110000",
    818 => "0101101110100000",
    819 => "0101111000000000",
    820 => "0110000001110000",
    821 => "0110001011100000",
    822 => "0110010101010000",
    823 => "0110011111010000",
    824 => "0110101001000000",
    825 => "0110110011000000",
    826 => "0110111101000000",
    827 => "0111000111000000",
    828 => "0111010001000000",
    829 => "0111011011000000",
    830 => "0111100101000000",
    831 => "0111101111000000",
    832 => "0111111001000000",
    833 => "1000000011010000",
    834 => "1000001101010000",
    835 => "1000010111010000",
    836 => "1000100001010000",
    837 => "1000101011010000",
    838 => "1000110101010000",
    839 => "1000111111010000",
    840 => "1001001001010000",
    841 => "1001010011010000",
    842 => "1001011101000000",
    843 => "1001100111000000",
    844 => "1001110000110000",
    845 => "1001111010100000",
    846 => "1010000100010000",
    847 => "1010001110000000",
    848 => "1010010111100000",
    849 => "1010100001010000",
    850 => "1010101010110000",
    851 => "1010110100000000",
    852 => "1010111101100000",
    853 => "1011000110110000",
    854 => "1011010000000000",
    855 => "1011011001010000",
    856 => "1011100010010000",
    857 => "1011101011010000",
    858 => "1011110100000000",
    859 => "1011111100110000",
    860 => "1100000101100000",
    861 => "1100001110000000",
    862 => "1100010110100000",
    863 => "1100011111000000",
    864 => "1100100111010000",
    865 => "1100101111100000",
    866 => "1100110111100000",
    867 => "1100111111010000",
    868 => "1101000111000000",
    869 => "1101001110110000",
    870 => "1101010110010000",
    871 => "1101011101110000",
    872 => "1101100101000000",
    873 => "1101101100010000",
    874 => "1101110011000000",
    875 => "1101111010000000",
    876 => "1110000000110000",
    877 => "1110000111010000",
    878 => "1110001101110000",
    879 => "1110010011110000",
    880 => "1110011010000000",
    881 => "1110100000000000",
    882 => "1110100101110000",
    883 => "1110101011010000",
    884 => "1110110000110000",
    885 => "1110110110000000",
    886 => "1110111011010000",
    887 => "1111000000000000",
    888 => "1111000100110000",
    889 => "1111001001100000",
    890 => "1111001101110000",
    891 => "1111010010000000",
    892 => "1111010110010000",
    893 => "1111011010000000",
    894 => "1111011101110000",
    895 => "1111100001010000",
    896 => "1111100100100000",
    897 => "1111100111110000",
    898 => "1111101010110000",
    899 => "1111101101100000",
    900 => "1111110000000000",
    901 => "1111110010010000",
    902 => "1111110100100000",
    903 => "1111110110100000",
    904 => "1111111000010000",
    905 => "1111111010000000",
    906 => "1111111011010000",
    907 => "1111111100100000",
    908 => "1111111101100000",
    909 => "1111111110100000",
    910 => "1111111111000000",
    911 => "1111111111100000",
    912 => "1111111111110000",
    913 => "1111111111110000",
    914 => "1111111111100000",
    915 => "1111111111010000",
    916 => "1111111110110000",
    917 => "1111111110000000",
    918 => "1111111101000000",
    919 => "1111111011110000",
    920 => "1111111010100000",
    921 => "1111111001000000",
    922 => "1111110111010000",
    923 => "1111110101010000",
    924 => "1111110011010000",
    925 => "1111110000110000",
    926 => "1111101110010000",
    927 => "1111101011110000",
    928 => "1111101000110000",
    929 => "1111100101110000",
    930 => "1111100010100000",
    931 => "1111011111000000",
    932 => "1111011011010000",
    933 => "1111010111100000",
    934 => "1111010011100000",
    935 => "1111001111010000",
    936 => "1111001011000000",
    937 => "1111000110100000",
    938 => "1111000001110000",
    939 => "1110111101000000",
    940 => "1110110111110000",
    941 => "1110110010100000",
    942 => "1110101101010000",
    943 => "1110100111110000",
    944 => "1110100010000000",
    945 => "1110011100000000",
    946 => "1110010110000000",
    947 => "1110001111110000",
    948 => "1110001001100000",
    949 => "1110000011000000",
    950 => "1101111100010000",
    951 => "1101110101100000",
    952 => "1101101110100000",
    953 => "1101100111100000",
    954 => "1101100000010000",
    955 => "1101011001000000",
    956 => "1101010001100000",
    957 => "1101001001110000",
    958 => "1101000010000000",
    959 => "1100111010010000",
    960 => "1100110010010000",
    961 => "1100101010000000",
    962 => "1100100010000000",
    963 => "1100011001100000",
    964 => "1100010001000000",
    965 => "1100001000100000",
    966 => "1100000000000000",
    967 => "1011110111010000",
    968 => "1011101110010000",
    969 => "1011100101010000",
    970 => "1011011100010000",
    971 => "1011010011010000",
    972 => "1011001010000000",
    973 => "1011000000110000",
    974 => "1010110111100000",
    975 => "1010101110000000",
    976 => "1010100100100000",
    977 => "1010011011000000",
    978 => "1010010001010000",
    979 => "1010000111110000",
    980 => "1001111110000000",
    981 => "1001110100010000",
    982 => "1001101010100000",
    983 => "1001100000100000",
    984 => "1001010110110000",
    985 => "1001001100110000",
    986 => "1001000010110000",
    987 => "1000111000110000",
    988 => "1000101110110000",
    989 => "1000100100110000",
    990 => "1000011010110000",
    991 => "1000010000110000",
    992 => "1000000110110000",
    993 => "0111111100100000",
    994 => "0111110010100000",
    995 => "0111101000100000",
    996 => "0111011110100000",
    997 => "0111010100100000",
    998 => "0111001010100000",
    999 => "0111000000100000",
    1000 => "0110110110100000",
    1001 => "0110101100100000",
    1002 => "0110100010110000",
    1003 => "0110011000110000",
    1004 => "0110001111000000",
    1005 => "0110000101010000",
    1006 => "0101111011100000",
    1007 => "0101110001110000",
    1008 => "0101101000010000",
    1009 => "0101011110100000",
    1010 => "0101010101000000",
    1011 => "0101001011110000",
    1012 => "0101000010010000",
    1013 => "0100111001000000",
    1014 => "0100101111110000",
    1015 => "0100100110100000",
    1016 => "0100011101100000",
    1017 => "0100010100100000",
    1018 => "0100001011110000",
    1019 => "0100000011000000",
    1020 => "0011111010010000",
    1021 => "0011110001110000",
    1022 => "0011101001010000",
    1023 => "0011100000110000",
    1024 => "0011011000100000",
    1025 => "0011010000010000",
    1026 => "0011001000010000",
    1027 => "0011000000100000",
    1028 => "0010111000110000",
    1029 => "0010110001000000",
    1030 => "0010101001100000",
    1031 => "0010100010000000",
    1032 => "0010011010110000",
    1033 => "0010010011100000",
    1034 => "0010001100110000",
    1035 => "0010000101110000",
    1036 => "0001111111000000",
    1037 => "0001111000100000",
    1038 => "0001110010000000",
    1039 => "0001101100000000",
    1040 => "0001100101110000",
    1041 => "0001011111110000",
    1042 => "0001011010000000",
    1043 => "0001010100100000",
    1044 => "0001001111000000",
    1045 => "0001001001110000",
    1046 => "0001000100100000",
    1047 => "0000111111110000",
    1048 => "0000111011000000",
    1049 => "0000110110010000",
    1050 => "0000110010000000",
    1051 => "0000101101110000",
    1052 => "0000101001100000",
    1053 => "0000100101110000",
    1054 => "0000100010000000",
    1055 => "0000011110100000",
    1056 => "0000011011010000",
    1057 => "0000011000000000",
    1058 => "0000010101000000",
    1059 => "0000010010010000",
    1060 => "0000001111110000",
    1061 => "0000001101100000",
    1062 => "0000001011010000",
    1063 => "0000001001010000",
    1064 => "0000000111100000",
    1065 => "0000000101110000",
    1066 => "0000000100100000",
    1067 => "0000000011010000",
    1068 => "0000000010010000",
    1069 => "0000000001010000",
    1070 => "0000000000110000",
    1071 => "0000000000010000",
    1072 => "0000000000000000",
    1073 => "0000000000000000",
    1074 => "0000000000010000",
    1075 => "0000000000100000",
    1076 => "0000000001000000",
    1077 => "0000000001110000",
    1078 => "0000000010110000",
    1079 => "0000000100000000",
    1080 => "0000000101010000",
    1081 => "0000000110110000",
    1082 => "0000001000100000",
    1083 => "0000001010100000",
    1084 => "0000001100100000",
    1085 => "0000001111000000",
    1086 => "0000010001100000",
    1087 => "0000010100000000",
    1088 => "0000010111000000",
    1089 => "0000011010000000",
    1090 => "0000011101010000",
    1091 => "0000100000110000",
    1092 => "0000100100100000",
    1093 => "0000101000010000",
    1094 => "0000101100010000",
    1095 => "0000110000100000",
    1096 => "0000110100110000",
    1097 => "0000111001010000",
    1098 => "0000111110000000",
    1099 => "0001000010110000",
    1100 => "0001001000000000",
    1101 => "0001001101010000",
    1102 => "0001010010100000",
    1103 => "0001011000000000",
    1104 => "0001011101110000",
    1105 => "0001100011110000",
    1106 => "0001101001110000",
    1107 => "0001110000000000",
    1108 => "0001110110010000",
    1109 => "0001111100110000",
    1110 => "0010000011100000",
    1111 => "0010001010010000",
    1112 => "0010010001010000",
    1113 => "0010011000010000",
    1114 => "0010011111100000",
    1115 => "0010100110110000",
    1116 => "0010101110010000",
    1117 => "0010110110000000",
    1118 => "0010111101110000",
    1119 => "0011000101100000",
    1120 => "0011001101100000",
    1121 => "0011010101110000",
    1122 => "0011011101110000",
    1123 => "0011100110010000",
    1124 => "0011101110110000",
    1125 => "0011110111010000",
    1126 => "0011111111110000",
    1127 => "0100001000100000",
    1128 => "0100010001100000",
    1129 => "0100011010100000",
    1130 => "0100100011100000",
    1131 => "0100101100100000",
    1132 => "0100110101110000",
    1133 => "0100111111000000",
    1134 => "0101001000010000",
    1135 => "0101010001110000",
    1136 => "0101011011010000",
    1137 => "0101100100110000",
    1138 => "0101101110100000",
    1139 => "0101111000000000",
    1140 => "0110000001110000",
    1141 => "0110001011100000",
    1142 => "0110010101010000",
    1143 => "0110011111010000",
    1144 => "0110101001000000",
    1145 => "0110110011000000",
    1146 => "0110111101000000",
    1147 => "0111000111000000",
    1148 => "0111010001000000",
    1149 => "0111011011000000",
    1150 => "0111100101000000",
    1151 => "0111101111000000",
    1152 => "0111111001000000",
    1153 => "1000000011010000",
    1154 => "1000001101010000",
    1155 => "1000010111010000",
    1156 => "1000100001010000",
    1157 => "1000101011010000",
    1158 => "1000110101010000",
    1159 => "1000111111010000",
    1160 => "1001001001010000",
    1161 => "1001010011010000",
    1162 => "1001011101000000",
    1163 => "1001100111000000",
    1164 => "1001110000110000",
    1165 => "1001111010100000",
    1166 => "1010000100010000",
    1167 => "1010001110000000",
    1168 => "1010010111100000",
    1169 => "1010100001010000",
    1170 => "1010101010110000",
    1171 => "1010110100000000",
    1172 => "1010111101100000",
    1173 => "1011000110110000",
    1174 => "1011010000000000",
    1175 => "1011011001010000",
    1176 => "1011100010010000",
    1177 => "1011101011010000",
    1178 => "1011110100000000",
    1179 => "1011111100110000",
    1180 => "1100000101100000",
    1181 => "1100001110000000",
    1182 => "1100010110100000",
    1183 => "1100011111000000",
    1184 => "1100100111010000",
    1185 => "1100101111100000",
    1186 => "1100110111100000",
    1187 => "1100111111010000",
    1188 => "1101000111000000",
    1189 => "1101001110110000",
    1190 => "1101010110010000",
    1191 => "1101011101110000",
    1192 => "1101100101000000",
    1193 => "1101101100010000",
    1194 => "1101110011000000",
    1195 => "1101111010000000",
    1196 => "1110000000110000",
    1197 => "1110000111010000",
    1198 => "1110001101110000",
    1199 => "1110010011110000",
    1200 => "1110011010000000",
    1201 => "1110100000000000",
    1202 => "1110100101110000",
    1203 => "1110101011010000",
    1204 => "1110110000110000",
    1205 => "1110110110000000",
    1206 => "1110111011010000",
    1207 => "1111000000000000",
    1208 => "1111000100110000",
    1209 => "1111001001100000",
    1210 => "1111001101110000",
    1211 => "1111010010000000",
    1212 => "1111010110010000",
    1213 => "1111011010000000",
    1214 => "1111011101110000",
    1215 => "1111100001010000",
    1216 => "1111100100100000",
    1217 => "1111100111110000",
    1218 => "1111101010110000",
    1219 => "1111101101100000",
    1220 => "1111110000000000",
    1221 => "1111110010010000",
    1222 => "1111110100100000",
    1223 => "1111110110100000",
    1224 => "1111111000010000",
    1225 => "1111111010000000",
    1226 => "1111111011010000",
    1227 => "1111111100100000",
    1228 => "1111111101100000",
    1229 => "1111111110100000",
    1230 => "1111111111000000",
    1231 => "1111111111100000",
    1232 => "1111111111110000",
    1233 => "1111111111110000",
    1234 => "1111111111100000",
    1235 => "1111111111010000",
    1236 => "1111111110110000",
    1237 => "1111111110000000",
    1238 => "1111111101000000",
    1239 => "1111111011110000",
    1240 => "1111111010100000",
    1241 => "1111111001000000",
    1242 => "1111110111010000",
    1243 => "1111110101010000",
    1244 => "1111110011010000",
    1245 => "1111110000110000",
    1246 => "1111101110010000",
    1247 => "1111101011110000",
    1248 => "1111101000110000",
    1249 => "1111100101110000",
    1250 => "1111100010100000",
    1251 => "1111011111000000",
    1252 => "1111011011010000",
    1253 => "1111010111100000",
    1254 => "1111010011100000",
    1255 => "1111001111010000",
    1256 => "1111001011000000",
    1257 => "1111000110100000",
    1258 => "1111000001110000",
    1259 => "1110111101000000",
    1260 => "1110110111110000",
    1261 => "1110110010100000",
    1262 => "1110101101010000",
    1263 => "1110100111110000",
    1264 => "1110100010000000",
    1265 => "1110011100000000",
    1266 => "1110010110000000",
    1267 => "1110001111110000",
    1268 => "1110001001100000",
    1269 => "1110000011000000",
    1270 => "1101111100010000",
    1271 => "1101110101100000",
    1272 => "1101101110100000",
    1273 => "1101100111100000",
    1274 => "1101100000010000",
    1275 => "1101011001000000",
    1276 => "1101010001100000",
    1277 => "1101001001110000",
    1278 => "1101000010000000",
    1279 => "1100111010010000",
    1280 => "1100110010010000",
    1281 => "1100101010000000",
    1282 => "1100100010000000",
    1283 => "1100011001100000",
    1284 => "1100010001000000",
    1285 => "1100001000100000",
    1286 => "1100000000000000",
    1287 => "1011110111010000",
    1288 => "1011101110010000",
    1289 => "1011100101010000",
    1290 => "1011011100010000",
    1291 => "1011010011010000",
    1292 => "1011001010000000",
    1293 => "1011000000110000",
    1294 => "1010110111100000",
    1295 => "1010101110000000",
    1296 => "1010100100100000",
    1297 => "1010011011000000",
    1298 => "1010010001010000",
    1299 => "1010000111110000",
    1300 => "1001111110000000",
    1301 => "1001110100010000",
    1302 => "1001101010100000",
    1303 => "1001100000100000",
    1304 => "1001010110110000",
    1305 => "1001001100110000",
    1306 => "1001000010110000",
    1307 => "1000111000110000",
    1308 => "1000101110110000",
    1309 => "1000100100110000",
    1310 => "1000011010110000",
    1311 => "1000010000110000",
    1312 => "1000000110110000",
    1313 => "0111111100100000",
    1314 => "0111110010100000",
    1315 => "0111101000100000",
    1316 => "0111011110100000",
    1317 => "0111010100100000",
    1318 => "0111001010100000",
    1319 => "0111000000100000",
    1320 => "0110110110100000",
    1321 => "0110101100100000",
    1322 => "0110100010110000",
    1323 => "0110011000110000",
    1324 => "0110001111000000",
    1325 => "0110000101010000",
    1326 => "0101111011100000",
    1327 => "0101110001110000",
    1328 => "0101101000010000",
    1329 => "0101011110100000",
    1330 => "0101010101000000",
    1331 => "0101001011110000",
    1332 => "0101000010010000",
    1333 => "0100111001000000",
    1334 => "0100101111110000",
    1335 => "0100100110100000",
    1336 => "0100011101100000",
    1337 => "0100010100100000",
    1338 => "0100001011110000",
    1339 => "0100000011000000",
    1340 => "0011111010010000",
    1341 => "0011110001110000",
    1342 => "0011101001010000",
    1343 => "0011100000110000",
    1344 => "0011011000100000",
    1345 => "0011010000010000",
    1346 => "0011001000010000",
    1347 => "0011000000100000",
    1348 => "0010111000110000",
    1349 => "0010110001000000",
    1350 => "0010101001100000",
    1351 => "0010100010000000",
    1352 => "0010011010110000",
    1353 => "0010010011100000",
    1354 => "0010001100110000",
    1355 => "0010000101110000",
    1356 => "0001111111000000",
    1357 => "0001111000100000",
    1358 => "0001110010000000",
    1359 => "0001101100000000",
    1360 => "0001100101110000",
    1361 => "0001011111110000",
    1362 => "0001011010000000",
    1363 => "0001010100100000",
    1364 => "0001001111000000",
    1365 => "0001001001110000",
    1366 => "0001000100100000",
    1367 => "0000111111110000",
    1368 => "0000111011000000",
    1369 => "0000110110010000",
    1370 => "0000110010000000",
    1371 => "0000101101110000",
    1372 => "0000101001100000",
    1373 => "0000100101110000",
    1374 => "0000100010000000",
    1375 => "0000011110100000",
    1376 => "0000011011010000",
    1377 => "0000011000000000",
    1378 => "0000010101000000",
    1379 => "0000010010010000",
    1380 => "0000001111110000",
    1381 => "0000001101100000",
    1382 => "0000001011010000",
    1383 => "0000001001010000",
    1384 => "0000000111100000",
    1385 => "0000000101110000",
    1386 => "0000000100100000",
    1387 => "0000000011010000",
    1388 => "0000000010010000",
    1389 => "0000000001010000",
    1390 => "0000000000110000",
    1391 => "0000000000010000",
    1392 => "0000000000000000",
    1393 => "0000000000000000",
    1394 => "0000000000010000",
    1395 => "0000000000100000",
    1396 => "0000000001000000",
    1397 => "0000000001110000",
    1398 => "0000000010110000",
    1399 => "0000000100000000",
    1400 => "0000000101010000",
    1401 => "0000000110110000",
    1402 => "0000001000100000",
    1403 => "0000001010100000",
    1404 => "0000001100100000",
    1405 => "0000001111000000",
    1406 => "0000010001100000",
    1407 => "0000010100000000",
    1408 => "0000010111000000",
    1409 => "0000011010000000",
    1410 => "0000011101010000",
    1411 => "0000100000110000",
    1412 => "0000100100100000",
    1413 => "0000101000010000",
    1414 => "0000101100010000",
    1415 => "0000110000100000",
    1416 => "0000110100110000",
    1417 => "0000111001010000",
    1418 => "0000111110000000",
    1419 => "0001000010110000",
    1420 => "0001001000000000",
    1421 => "0001001101010000",
    1422 => "0001010010100000",
    1423 => "0001011000000000",
    1424 => "0001011101110000",
    1425 => "0001100011110000",
    1426 => "0001101001110000",
    1427 => "0001110000000000",
    1428 => "0001110110010000",
    1429 => "0001111100110000",
    1430 => "0010000011100000",
    1431 => "0010001010010000",
    1432 => "0010010001010000",
    1433 => "0010011000010000",
    1434 => "0010011111100000",
    1435 => "0010100110110000",
    1436 => "0010101110010000",
    1437 => "0010110110000000",
    1438 => "0010111101110000",
    1439 => "0011000101100000",
    1440 => "0011001101100000",
    1441 => "0011010101110000",
    1442 => "0011011101110000",
    1443 => "0011100110010000",
    1444 => "0011101110110000",
    1445 => "0011110111010000",
    1446 => "0011111111110000",
    1447 => "0100001000100000",
    1448 => "0100010001100000",
    1449 => "0100011010100000",
    1450 => "0100100011100000",
    1451 => "0100101100100000",
    1452 => "0100110101110000",
    1453 => "0100111111000000",
    1454 => "0101001000010000",
    1455 => "0101010001110000",
    1456 => "0101011011010000",
    1457 => "0101100100110000",
    1458 => "0101101110100000",
    1459 => "0101111000000000",
    1460 => "0110000001110000",
    1461 => "0110001011100000",
    1462 => "0110010101010000",
    1463 => "0110011111010000",
    1464 => "0110101001000000",
    1465 => "0110110011000000",
    1466 => "0110111101000000",
    1467 => "0111000111000000",
    1468 => "0111010001000000",
    1469 => "0111011011000000",
    1470 => "0111100101000000",
    1471 => "0111101111000000",
    1472 => "0111111001000000",
    1473 => "1000000011010000",
    1474 => "1000001101010000",
    1475 => "1000010111010000",
    1476 => "1000100001010000",
    1477 => "1000101011010000",
    1478 => "1000110101010000",
    1479 => "1000111111010000",
    1480 => "1001001001010000",
    1481 => "1001010011010000",
    1482 => "1001011101000000",
    1483 => "1001100111000000",
    1484 => "1001110000110000",
    1485 => "1001111010100000",
    1486 => "1010000100010000",
    1487 => "1010001110000000",
    1488 => "1010010111100000",
    1489 => "1010100001010000",
    1490 => "1010101010110000",
    1491 => "1010110100000000",
    1492 => "1010111101100000",
    1493 => "1011000110110000",
    1494 => "1011010000000000",
    1495 => "1011011001010000",
    1496 => "1011100010010000",
    1497 => "1011101011010000",
    1498 => "1011110100000000",
    1499 => "1011111100110000",
    1500 => "1100000101100000",
    1501 => "1100001110000000",
    1502 => "1100010110100000",
    1503 => "1100011111000000",
    1504 => "1100100111010000",
    1505 => "1100101111100000",
    1506 => "1100110111100000",
    1507 => "1100111111010000",
    1508 => "1101000111000000",
    1509 => "1101001110110000",
    1510 => "1101010110010000",
    1511 => "1101011101110000",
    1512 => "1101100101000000",
    1513 => "1101101100010000",
    1514 => "1101110011000000",
    1515 => "1101111010000000",
    1516 => "1110000000110000",
    1517 => "1110000111010000",
    1518 => "1110001101110000",
    1519 => "1110010011110000",
    1520 => "1110011010000000",
    1521 => "1110100000000000",
    1522 => "1110100101110000",
    1523 => "1110101011010000",
    1524 => "1110110000110000",
    1525 => "1110110110000000",
    1526 => "1110111011010000",
    1527 => "1111000000000000",
    1528 => "1111000100110000",
    1529 => "1111001001100000",
    1530 => "1111001101110000",
    1531 => "1111010010000000",
    1532 => "1111010110010000",
    1533 => "1111011010000000",
    1534 => "1111011101110000",
    1535 => "1111100001010000",
    1536 => "1111100100100000",
    1537 => "1111100111110000",
    1538 => "1111101010110000",
    1539 => "1111101101100000",
    1540 => "1111110000000000",
    1541 => "1111110010010000",
    1542 => "1111110100100000",
    1543 => "1111110110100000",
    1544 => "1111111000010000",
    1545 => "1111111010000000",
    1546 => "1111111011010000",
    1547 => "1111111100100000",
    1548 => "1111111101100000",
    1549 => "1111111110100000",
    1550 => "1111111111000000",
    1551 => "1111111111100000",
    1552 => "1111111111110000",
    1553 => "1111111111110000",
    1554 => "1111111111100000",
    1555 => "1111111111010000",
    1556 => "1111111110110000",
    1557 => "1111111110000000",
    1558 => "1111111101000000",
    1559 => "1111111011110000",
    1560 => "1111111010100000",
    1561 => "1111111001000000",
    1562 => "1111110111010000",
    1563 => "1111110101010000",
    1564 => "1111110011010000",
    1565 => "1111110000110000",
    1566 => "1111101110010000",
    1567 => "1111101011110000",
    1568 => "1111101000110000",
    1569 => "1111100101110000",
    1570 => "1111100010100000",
    1571 => "1111011111000000",
    1572 => "1111011011010000",
    1573 => "1111010111100000",
    1574 => "1111010011100000",
    1575 => "1111001111010000",
    1576 => "1111001011000000",
    1577 => "1111000110100000",
    1578 => "1111000001110000",
    1579 => "1110111101000000",
    1580 => "1110110111110000",
    1581 => "1110110010100000",
    1582 => "1110101101010000",
    1583 => "1110100111110000",
    1584 => "1110100010000000",
    1585 => "1110011100000000",
    1586 => "1110010110000000",
    1587 => "1110001111110000",
    1588 => "1110001001100000",
    1589 => "1110000011000000",
    1590 => "1101111100010000",
    1591 => "1101110101100000",
    1592 => "1101101110100000",
    1593 => "1101100111100000",
    1594 => "1101100000010000",
    1595 => "1101011001000000",
    1596 => "1101010001100000",
    1597 => "1101001001110000",
    1598 => "1101000010000000",
    1599 => "1100111010010000"
    );
BEGIN
    PROCESS (clk)
    BEGIN
        IF rising_edge(clk) THEN
            data_out <= rom(address);
        END IF;
    END PROCESS;
END beh;